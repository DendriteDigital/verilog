module CharSet(
	input		wire				clock,
	input		wire	[ 7:0]	char,
	output	reg	[31:0]	pixels
);
	
	initial begin
		pixels<=32'd0;
	end
	
	always@(posedge clock)begin
		pixels<=rom[char];
	end
	
	wire[31:0]rom[255:0];

assign rom[  0]={8'b00000000,
                 8'b00110110,
                 8'b01111111,
                 8'b01111111};
assign rom[  1]={8'b00111110,
                 8'b00011100,
                 8'b00001000,
                 8'b00000000};

assign rom[  2]={8'b00011000,
                 8'b00011000,
                 8'b00011000,
                 8'b00011111};
assign rom[  3]={8'b00011111,
                 8'b00011000,
                 8'b00011000,
                 8'b00011000};

assign rom[  4]={8'b00000011,
                 8'b00000011,
                 8'b00000011,
                 8'b00000011};
assign rom[  5]={8'b00000011,
                 8'b00000011,
                 8'b00000011,
                 8'b00000011};

assign rom[  6]={8'b00011000,
                 8'b00011000,
                 8'b00011000,
                 8'b11111000};
assign rom[  7]={8'b11111000,
                 8'b00000000,
                 8'b00000000,
                 8'b00000000};

assign rom[  8]={8'b00011000,
                 8'b00011000,
                 8'b00011000,
                 8'b11111000};
assign rom[  9]={8'b11111000,
                 8'b00011000,
                 8'b00011000,
                 8'b00011000};

assign rom[ 10]={8'b00000000,
                 8'b00000000,
                 8'b00000000,
                 8'b11111000};
assign rom[ 11]={8'b11111000,
                 8'b00011000,
                 8'b00011000,
                 8'b00011000};

assign rom[ 12]={8'b00000011,
                 8'b00000111,
                 8'b00001110,
                 8'b00011100};
assign rom[ 13]={8'b00111000,
                 8'b01110000,
                 8'b11100000,
                 8'b11000000};

assign rom[ 14]={8'b11000000,
                 8'b11100000,
                 8'b01110000,
                 8'b00111000};
assign rom[ 15]={8'b00011100,
                 8'b00001110,
                 8'b00000111,
                 8'b00000011};

assign rom[ 16]={8'b00000001,
                 8'b00000011,
                 8'b00000111,
                 8'b00001111};
assign rom[ 17]={8'b00011111,
                 8'b00111111,
                 8'b01111111,
                 8'b11111111};

assign rom[ 18]={8'b00000000,
                 8'b00000000,
                 8'b00000000,
                 8'b00000000};
assign rom[ 19]={8'b00001111,
                 8'b00001111,
                 8'b00001111,
                 8'b00001111};

assign rom[ 20]={8'b10000000,
                 8'b11000000,
                 8'b11100000,
                 8'b11110000};
assign rom[ 21]={8'b11111000,
                 8'b11111100,
                 8'b11111110,
                 8'b11111111};

assign rom[ 22]={8'b00001111,
                 8'b00001111,
                 8'b00001111,
                 8'b00001111};
assign rom[ 23]={8'b00000000,
                 8'b00000000,
                 8'b00000000,
                 8'b00000000};

assign rom[ 24]={8'b11110000,
                 8'b11110000,
                 8'b11110000,
                 8'b11110000};
assign rom[ 25]={8'b00000000,
                 8'b00000000,
                 8'b00000000,
                 8'b00000000};

assign rom[ 26]={8'b11111111,
                 8'b11111111,
                 8'b00000000,
                 8'b00000000};
assign rom[ 27]={8'b00000000,
                 8'b00000000,
                 8'b00000000,
                 8'b00000000};

assign rom[ 28]={8'b00000000,
                 8'b00000000,
                 8'b00000000,
                 8'b00000000};
assign rom[ 29]={8'b00000000,
                 8'b00000000,
                 8'b11111111,
                 8'b11111111};

assign rom[ 30]={8'b00000000,
                 8'b00000000,
                 8'b00000000,
                 8'b00000000};
assign rom[ 31]={8'b11110000,
                 8'b11110000,
                 8'b11110000,
                 8'b11110000};

assign rom[ 32]={8'b00000000,
                 8'b00011100,
                 8'b00011100,
                 8'b01110111};
assign rom[ 33]={8'b01110111,
                 8'b00001000,
                 8'b00011100,
                 8'b00000000};

assign rom[ 34]={8'b00000000,
                 8'b00000000,
                 8'b00000000,
                 8'b00011111};
assign rom[ 35]={8'b00011111,
                 8'b00011000,
                 8'b00011000,
                 8'b00011000};

assign rom[ 36]={8'b00000000,
                 8'b00000000,
                 8'b00000000,
                 8'b11111111};
assign rom[ 37]={8'b11111111,
                 8'b00000000,
                 8'b00000000,
                 8'b00000000};

assign rom[ 38]={8'b00011000,
                 8'b00011000,
                 8'b00011000,
                 8'b11111111};
assign rom[ 39]={8'b11111111,
                 8'b00011000,
                 8'b00011000,
                 8'b00011000};

assign rom[ 40]={8'b00000000,
                 8'b00000000,
                 8'b00111100,
                 8'b01111110};
assign rom[ 41]={8'b01111110,
                 8'b01111110,
                 8'b00111100,
                 8'b00000000};

assign rom[ 42]={8'b00000000,
                 8'b00000000,
                 8'b00000000,
                 8'b00000000};
assign rom[ 43]={8'b11111111,
                 8'b11111111,
                 8'b11111111,
                 8'b11111111};

assign rom[ 44]={8'b11000000,
                 8'b11000000,
                 8'b11000000,
                 8'b11000000};
assign rom[ 45]={8'b11000000,
                 8'b11000000,
                 8'b11000000,
                 8'b11000000};

assign rom[ 46]={8'b00000000,
                 8'b00000000,
                 8'b00000000,
                 8'b11111111};
assign rom[ 47]={8'b11111111,
                 8'b00011000,
                 8'b00011000,
                 8'b00011000};

assign rom[ 48]={8'b00011000,
                 8'b00011000,
                 8'b00011000,
                 8'b11111111};
assign rom[ 49]={8'b11111111,
                 8'b00000000,
                 8'b00000000,
                 8'b00000000};

assign rom[ 50]={8'b11110000,
                 8'b11110000,
                 8'b11110000,
                 8'b11110000};
assign rom[ 51]={8'b11110000,
                 8'b11110000,
                 8'b11110000,
                 8'b11110000};

assign rom[ 52]={8'b00011000,
                 8'b00011000,
                 8'b00011000,
                 8'b00011111};
assign rom[ 53]={8'b00011111,
                 8'b00000000,
                 8'b00000000,
                 8'b00000000};

assign rom[ 54]={8'b01111000,
                 8'b01100000,
                 8'b01111000,
                 8'b01100000};
assign rom[ 55]={8'b01111110,
                 8'b00011000,
                 8'b00011110,
                 8'b00000000};

assign rom[ 56]={8'b00000000,
                 8'b00011000,
                 8'b00111100,
                 8'b01111110};
assign rom[ 57]={8'b00011000,
                 8'b00011000,
                 8'b00011000,
                 8'b00000000};

assign rom[ 58]={8'b00000000,
                 8'b00011000,
                 8'b00011000,
                 8'b00011000};
assign rom[ 59]={8'b01111110,
                 8'b00111100,
                 8'b00011000,
                 8'b00000000};

assign rom[ 60]={8'b00000000,
                 8'b00011000,
                 8'b00110000,
                 8'b01111110};
assign rom[ 61]={8'b00110000,
                 8'b00011000,
                 8'b00000000,
                 8'b00000000};

assign rom[ 62]={8'b00000000,
                 8'b00011000,
                 8'b00001100,
                 8'b01111110};
assign rom[ 63]={8'b00001100,
                 8'b00011000,
                 8'b00000000,
                 8'b00000000};

assign rom[ 64]={8'b00000000,
                 8'b00000000,
                 8'b00000000,
                 8'b00000000};
assign rom[ 65]={8'b00000000,
                 8'b00000000,
                 8'b00000000,
                 8'b00000000};

assign rom[ 66]={8'b00000000,
                 8'b00011000,
                 8'b00011000,
                 8'b00011000};
assign rom[ 67]={8'b00011000,
                 8'b00000000,
                 8'b00011000,
                 8'b00000000};

assign rom[ 68]={8'b00000000,
                 8'b01100110,
                 8'b01100110,
                 8'b01100110};
assign rom[ 69]={8'b00000000,
                 8'b00000000,
                 8'b00000000,
                 8'b00000000};

assign rom[ 70]={8'b00000000,
                 8'b01100110,
                 8'b11111111,
                 8'b01100110};
assign rom[ 71]={8'b01100110,
                 8'b11111111,
                 8'b01100110,
                 8'b00000000};

assign rom[ 72]={8'b00011000,
                 8'b00111110,
                 8'b01100000,
                 8'b00111100};
assign rom[ 73]={8'b00000110,
                 8'b01111100,
                 8'b00011000,
                 8'b00000000};

assign rom[ 74]={8'b00000000,
                 8'b01100110,
                 8'b01101100,
                 8'b00011000};
assign rom[ 75]={8'b00110000,
                 8'b01100110,
                 8'b01000110,
                 8'b00000000};

assign rom[ 76]={8'b00011100,
                 8'b00110110,
                 8'b00011100,
                 8'b00111000};
assign rom[ 77]={8'b01101111,
                 8'b01100110,
                 8'b00111011,
                 8'b00000000};

assign rom[ 78]={8'b00000000,
                 8'b00011000,
                 8'b00011000,
                 8'b00011000};
assign rom[ 79]={8'b00000000,
                 8'b00000000,
                 8'b00000000,
                 8'b00000000};

assign rom[ 80]={8'b00000000,
                 8'b00001110,
                 8'b00011100,
                 8'b00011000};
assign rom[ 81]={8'b00011000,
                 8'b00011100,
                 8'b00001110,
                 8'b00000000};

assign rom[ 82]={8'b00000000,
                 8'b01110000,
                 8'b00111000,
                 8'b00011000};
assign rom[ 83]={8'b00011000,
                 8'b00111000,
                 8'b01110000,
                 8'b00000000};

assign rom[ 84]={8'b00000000,
                 8'b01100110,
                 8'b00111100,
                 8'b11111111};
assign rom[ 85]={8'b00111100,
                 8'b01100110,
                 8'b00000000,
                 8'b00000000};

assign rom[ 86]={8'b00000000,
                 8'b00011000,
                 8'b00011000,
                 8'b01111110};
assign rom[ 87]={8'b00011000,
                 8'b00011000,
                 8'b00000000,
                 8'b00000000};

assign rom[ 88]={8'b00000000,
                 8'b00000000,
                 8'b00000000,
                 8'b00000000};
assign rom[ 89]={8'b00000000,
                 8'b00011000,
                 8'b00011000,
                 8'b00110000};

assign rom[ 90]={8'b00000000,
                 8'b00000000,
                 8'b00000000,
                 8'b01111110};
assign rom[ 91]={8'b00000000,
                 8'b00000000,
                 8'b00000000,
                 8'b00000000};

assign rom[ 92]={8'b00000000,
                 8'b00000000,
                 8'b00000000,
                 8'b00000000};
assign rom[ 93]={8'b00000000,
                 8'b00011000,
                 8'b00011000,
                 8'b00000000};

assign rom[ 94]={8'b00000000,
                 8'b00000110,
                 8'b00001100,
                 8'b00011000};
assign rom[ 95]={8'b00110000,
                 8'b01100000,
                 8'b01000000,
                 8'b00000000};

assign rom[ 96]={8'b00000000,
                 8'b00111100,
                 8'b01100110,
                 8'b01101110};
assign rom[ 97]={8'b01110110,
                 8'b01100110,
                 8'b00111100,
                 8'b00000000};

assign rom[ 98]={8'b00000000,
                 8'b00011000,
                 8'b00111000,
                 8'b00011000};
assign rom[ 99]={8'b00011000,
                 8'b00011000,
                 8'b01111110,
                 8'b00000000};

assign rom[100]={8'b00000000,
                 8'b00111100,
                 8'b01100110,
                 8'b00001100};
assign rom[101]={8'b00011000,
                 8'b00110000,
                 8'b01111110,
                 8'b00000000};

assign rom[102]={8'b00000000,
                 8'b01111110,
                 8'b00001100,
                 8'b00011000};
assign rom[103]={8'b00001100,
                 8'b01100110,
                 8'b00111100,
                 8'b00000000};

assign rom[104]={8'b00000000,
                 8'b00001100,
                 8'b00011100,
                 8'b00111100};
assign rom[105]={8'b01101100,
                 8'b01111110,
                 8'b00001100,
                 8'b00000000};

assign rom[106]={8'b00000000,
                 8'b01111110,
                 8'b01100000,
                 8'b01111100};
assign rom[107]={8'b00000110,
                 8'b01100110,
                 8'b00111100,
                 8'b00000000};

assign rom[108]={8'b00000000,
                 8'b00111100,
                 8'b01100000,
                 8'b01111100};
assign rom[109]={8'b01100110,
                 8'b01100110,
                 8'b00111100,
                 8'b00000000};

assign rom[110]={8'b00000000,
                 8'b01111110,
                 8'b00000110,
                 8'b00001100};
assign rom[111]={8'b00011000,
                 8'b00110000,
                 8'b00110000,
                 8'b00000000};

assign rom[112]={8'b00000000,
                 8'b00111100,
                 8'b01100110,
                 8'b00111100};
assign rom[113]={8'b01100110,
                 8'b01100110,
                 8'b00111100,
                 8'b00000000};

assign rom[114]={8'b00000000,
                 8'b00111100,
                 8'b01100110,
                 8'b00111110};
assign rom[115]={8'b00000110,
                 8'b00001100,
                 8'b00111000,
                 8'b00000000};

assign rom[116]={8'b00000000,
                 8'b00000000,
                 8'b00011000,
                 8'b00011000};
assign rom[117]={8'b00000000,
                 8'b00011000,
                 8'b00011000,
                 8'b00000000};

assign rom[118]={8'b00000000,
                 8'b00000000,
                 8'b00011000,
                 8'b00011000};
assign rom[119]={8'b00000000,
                 8'b00011000,
                 8'b00011000,
                 8'b00110000};

assign rom[120]={8'b00000110,
                 8'b00001100,
                 8'b00011000,
                 8'b00110000};
assign rom[121]={8'b00011000,
                 8'b00001100,
                 8'b00000110,
                 8'b00000000};

assign rom[122]={8'b00000000,
                 8'b00000000,
                 8'b01111110,
                 8'b00000000};
assign rom[123]={8'b00000000,
                 8'b01111110,
                 8'b00000000,
                 8'b00000000};

assign rom[124]={8'b01100000,
                 8'b00110000,
                 8'b00011000,
                 8'b00001100};
assign rom[125]={8'b00011000,
                 8'b00110000,
                 8'b01100000,
                 8'b00000000};

assign rom[126]={8'b00000000,
                 8'b00111100,
                 8'b01100110,
                 8'b00001100};
assign rom[127]={8'b00011000,
                 8'b00000000,
                 8'b00011000,
                 8'b00000000};

assign rom[128]={8'b00000000,
                 8'b00111100,
                 8'b01100110,
                 8'b01101110};
assign rom[129]={8'b01101110,
                 8'b01100000,
                 8'b00111110,
                 8'b00000000};

assign rom[130]={8'b00000000,
                 8'b00011000,
                 8'b00111100,
                 8'b01100110};
assign rom[131]={8'b01100110,
                 8'b01111110,
                 8'b01100110,
                 8'b00000000};

assign rom[132]={8'b00000000,
                 8'b01111100,
                 8'b01100110,
                 8'b01111100};
assign rom[133]={8'b01100110,
                 8'b01100110,
                 8'b01111100,
                 8'b00000000};

assign rom[134]={8'b00000000,
                 8'b00111100,
                 8'b01100110,
                 8'b01100000};
assign rom[135]={8'b01100000,
                 8'b01100110,
                 8'b00111100,
                 8'b00000000};

assign rom[136]={8'b00000000,
                 8'b01111000,
                 8'b01101100,
                 8'b01100110};
assign rom[137]={8'b01100110,
                 8'b01101100,
                 8'b01111000,
                 8'b00000000};

assign rom[138]={8'b00000000,
                 8'b01111110,
                 8'b01100000,
                 8'b01111100};
assign rom[139]={8'b01100000,
                 8'b01100000,
                 8'b01111110,
                 8'b00000000};

assign rom[140]={8'b00000000,
                 8'b01111110,
                 8'b01100000,
                 8'b01111100};
assign rom[141]={8'b01100000,
                 8'b01100000,
                 8'b01100000,
                 8'b00000000};

assign rom[142]={8'b00000000,
                 8'b00111110,
                 8'b01100000,
                 8'b01100000};
assign rom[143]={8'b01101110,
                 8'b01100110,
                 8'b00111110,
                 8'b00000000};

assign rom[144]={8'b00000000,
                 8'b01100110,
                 8'b01100110,
                 8'b01111110};
assign rom[145]={8'b01100110,
                 8'b01100110,
                 8'b01100110,
                 8'b00000000};

assign rom[146]={8'b00000000,
                 8'b01111110,
                 8'b00011000,
                 8'b00011000};
assign rom[147]={8'b00011000,
                 8'b00011000,
                 8'b01111110,
                 8'b00000000};

assign rom[148]={8'b00000000,
                 8'b00000110,
                 8'b00000110,
                 8'b00000110};
assign rom[149]={8'b00000110,
                 8'b01100110,
                 8'b00111100,
                 8'b00000000};

assign rom[150]={8'b00000000,
                 8'b01100110,
                 8'b01101100,
                 8'b01111000};
assign rom[151]={8'b01111000,
                 8'b01101100,
                 8'b01100110,
                 8'b00000000};

assign rom[152]={8'b00000000,
                 8'b01100000,
                 8'b01100000,
                 8'b01100000};
assign rom[153]={8'b01100000,
                 8'b01100000,
                 8'b01111110,
                 8'b00000000};

assign rom[154]={8'b00000000,
                 8'b01100011,
                 8'b01110111,
                 8'b01111111};
assign rom[155]={8'b01101011,
                 8'b01100011,
                 8'b01100011,
                 8'b00000000};

assign rom[156]={8'b00000000,
                 8'b01100110,
                 8'b01110110,
                 8'b01111110};
assign rom[157]={8'b01111110,
                 8'b01101110,
                 8'b01100110,
                 8'b00000000};

assign rom[158]={8'b00000000,
                 8'b00111100,
                 8'b01100110,
                 8'b01100110};
assign rom[159]={8'b01100110,
                 8'b01100110,
                 8'b00111100,
                 8'b00000000};

assign rom[160]={8'b00000000,
                 8'b01111100,
                 8'b01100110,
                 8'b01100110};
assign rom[161]={8'b01111100,
                 8'b01100000,
                 8'b01100000,
                 8'b00000000};

assign rom[162]={8'b00000000,
                 8'b00111100,
                 8'b01100110,
                 8'b01100110};
assign rom[163]={8'b01100110,
                 8'b01101100,
                 8'b00110110,
                 8'b00000000};

assign rom[164]={8'b00000000,
                 8'b01111100,
                 8'b01100110,
                 8'b01100110};
assign rom[165]={8'b01111100,
                 8'b01101100,
                 8'b01100110,
                 8'b00000000};

assign rom[166]={8'b00000000,
                 8'b00111100,
                 8'b01100000,
                 8'b00111100};
assign rom[167]={8'b00000110,
                 8'b00000110,
                 8'b00111100,
                 8'b00000000};

assign rom[168]={8'b00000000,
                 8'b01111110,
                 8'b00011000,
                 8'b00011000};
assign rom[169]={8'b00011000,
                 8'b00011000,
                 8'b00011000,
                 8'b00000000};

assign rom[170]={8'b00000000,
                 8'b01100110,
                 8'b01100110,
                 8'b01100110};
assign rom[171]={8'b01100110,
                 8'b01100110,
                 8'b01111110,
                 8'b00000000};

assign rom[172]={8'b00000000,
                 8'b01100110,
                 8'b01100110,
                 8'b01100110};
assign rom[173]={8'b01100110,
                 8'b00111100,
                 8'b00011000,
                 8'b00000000};

assign rom[174]={8'b00000000,
                 8'b01100011,
                 8'b01100011,
                 8'b01101011};
assign rom[175]={8'b01111111,
                 8'b01110111,
                 8'b01100011,
                 8'b00000000};

assign rom[176]={8'b00000000,
                 8'b01100110,
                 8'b01100110,
                 8'b00111100};
assign rom[177]={8'b00111100,
                 8'b01100110,
                 8'b01100110,
                 8'b00000000};

assign rom[178]={8'b00000000,
                 8'b01100110,
                 8'b01100110,
                 8'b00111100};
assign rom[179]={8'b00011000,
                 8'b00011000,
                 8'b00011000,
                 8'b00000000};

assign rom[180]={8'b00000000,
                 8'b01111110,
                 8'b00001100,
                 8'b00011000};
assign rom[181]={8'b00110000,
                 8'b01100000,
                 8'b01111110,
                 8'b00000000};

assign rom[182]={8'b00000000,
                 8'b00011110,
                 8'b00011000,
                 8'b00011000};
assign rom[183]={8'b00011000,
                 8'b00011000,
                 8'b00011110,
                 8'b00000000};

assign rom[184]={8'b00000000,
                 8'b01000000,
                 8'b01100000,
                 8'b00110000};
assign rom[185]={8'b00011000,
                 8'b00001100,
                 8'b00000110,
                 8'b00000000};

assign rom[186]={8'b00000000,
                 8'b01111000,
                 8'b00011000,
                 8'b00011000};
assign rom[187]={8'b00011000,
                 8'b00011000,
                 8'b01111000,
                 8'b00000000};

assign rom[188]={8'b00000000,
                 8'b00001000,
                 8'b00011100,
                 8'b00110110};
assign rom[189]={8'b01100011,
                 8'b00000000,
                 8'b00000000,
                 8'b00000000};

assign rom[190]={8'b00000000,
                 8'b00000000,
                 8'b00000000,
                 8'b00000000};
assign rom[191]={8'b00000000,
                 8'b00000000,
                 8'b11111111,
                 8'b00000000};

assign rom[192]={8'b00000000,
                 8'b00011000,
                 8'b00111100,
                 8'b01111110};
assign rom[193]={8'b01111110,
                 8'b00111100,
                 8'b00011000,
                 8'b00000000};

assign rom[194]={8'b00000000,
                 8'b00000000,
                 8'b00111100,
                 8'b00000110};
assign rom[195]={8'b00111110,
                 8'b01100110,
                 8'b00111110,
                 8'b00000000};

assign rom[196]={8'b00000000,
                 8'b01100000,
                 8'b01100000,
                 8'b01111100};
assign rom[197]={8'b01100110,
                 8'b01100110,
                 8'b01111100,
                 8'b00000000};

assign rom[198]={8'b00000000,
                 8'b00000000,
                 8'b00111100,
                 8'b01100000};
assign rom[199]={8'b01100000,
                 8'b01100000,
                 8'b00111100,
                 8'b00000000};

assign rom[200]={8'b00000000,
                 8'b00000110,
                 8'b00000110,
                 8'b00111110};
assign rom[201]={8'b01100110,
                 8'b01100110,
                 8'b00111110,
                 8'b00000000};

assign rom[202]={8'b00000000,
                 8'b00000000,
                 8'b00111100,
                 8'b01100110};
assign rom[203]={8'b01111110,
                 8'b01100000,
                 8'b00111100,
                 8'b00000000};

assign rom[204]={8'b00000000,
                 8'b00001110,
                 8'b00011000,
                 8'b00111110};
assign rom[205]={8'b00011000,
                 8'b00011000,
                 8'b00011000,
                 8'b00000000};

assign rom[206]={8'b00000000,
                 8'b00000000,
                 8'b00111110,
                 8'b01100110};
assign rom[207]={8'b01100110,
                 8'b00111110,
                 8'b00000110,
                 8'b01111100};

assign rom[208]={8'b00000000,
                 8'b01100000,
                 8'b01100000,
                 8'b01111100};
assign rom[209]={8'b01100110,
                 8'b01100110,
                 8'b01100110,
                 8'b00000000};

assign rom[210]={8'b00000000,
                 8'b00011000,
                 8'b00000000,
                 8'b00111000};
assign rom[211]={8'b00011000,
                 8'b00011000,
                 8'b00111100,
                 8'b00000000};

assign rom[212]={8'b00000000,
                 8'b00000110,
                 8'b00000000,
                 8'b00000110};
assign rom[213]={8'b00000110,
                 8'b00000110,
                 8'b00000110,
                 8'b00111100};

assign rom[214]={8'b00000000,
                 8'b01100000,
                 8'b01100000,
                 8'b01101100};
assign rom[215]={8'b01111000,
                 8'b01101100,
                 8'b01100110,
                 8'b00000000};

assign rom[216]={8'b00000000,
                 8'b00111000,
                 8'b00011000,
                 8'b00011000};
assign rom[217]={8'b00011000,
                 8'b00011000,
                 8'b00111100,
                 8'b00000000};

assign rom[218]={8'b00000000,
                 8'b00000000,
                 8'b01100110,
                 8'b01111111};
assign rom[219]={8'b01111111,
                 8'b01101011,
                 8'b01100011,
                 8'b00000000};

assign rom[220]={8'b00000000,
                 8'b00000000,
                 8'b01111100,
                 8'b01100110};
assign rom[221]={8'b01100110,
                 8'b01100110,
                 8'b01100110,
                 8'b00000000};

assign rom[222]={8'b00000000,
                 8'b00000000,
                 8'b00111100,
                 8'b01100110};
assign rom[223]={8'b01100110,
                 8'b01100110,
                 8'b00111100,
                 8'b00000000};

assign rom[224]={8'b00000000,
                 8'b00000000,
                 8'b01111100,
                 8'b01100110};
assign rom[225]={8'b01100110,
                 8'b01111100,
                 8'b01100000,
                 8'b01100000};

assign rom[226]={8'b00000000,
                 8'b00000000,
                 8'b00111110,
                 8'b01100110};
assign rom[227]={8'b01100110,
                 8'b00111110,
                 8'b00000110,
                 8'b00000110};

assign rom[228]={8'b00000000,
                 8'b00000000,
                 8'b01111100,
                 8'b01100110};
assign rom[229]={8'b01100000,
                 8'b01100000,
                 8'b01100000,
                 8'b00000000};

assign rom[230]={8'b00000000,
                 8'b00000000,
                 8'b00111110,
                 8'b01100000};
assign rom[231]={8'b00111100,
                 8'b00000110,
                 8'b01111100,
                 8'b00000000};

assign rom[232]={8'b00000000,
                 8'b00011000,
                 8'b01111110,
                 8'b00011000};
assign rom[233]={8'b00011000,
                 8'b00011000,
                 8'b00001110,
                 8'b00000000};

assign rom[234]={8'b00000000,
                 8'b00000000,
                 8'b01100110,
                 8'b01100110};
assign rom[235]={8'b01100110,
                 8'b01100110,
                 8'b00111110,
                 8'b00000000};

assign rom[236]={8'b00000000,
                 8'b00000000,
                 8'b01100110,
                 8'b01100110};
assign rom[237]={8'b01100110,
                 8'b00111100,
                 8'b00011000,
                 8'b00000000};

assign rom[238]={8'b00000000,
                 8'b00000000,
                 8'b01100011,
                 8'b01101011};
assign rom[239]={8'b01111111,
                 8'b00111110,
                 8'b00110110,
                 8'b00000000};

assign rom[240]={8'b00000000,
                 8'b00000000,
                 8'b01100110,
                 8'b00111100};
assign rom[241]={8'b00011000,
                 8'b00111100,
                 8'b01100110,
                 8'b00000000};

assign rom[242]={8'b00000000,
                 8'b00000000,
                 8'b01100110,
                 8'b01100110};
assign rom[243]={8'b01100110,
                 8'b00111110,
                 8'b00001100,
                 8'b01111000};

assign rom[244]={8'b00000000,
                 8'b00000000,
                 8'b01111110,
                 8'b00001100};
assign rom[245]={8'b00011000,
                 8'b00110000,
                 8'b01111110,
                 8'b00000000};

assign rom[246]={8'b00000000,
                 8'b00011000,
                 8'b00111100,
                 8'b01111110};
assign rom[247]={8'b01111110,
                 8'b00011000,
                 8'b00111100,
                 8'b00000000};

assign rom[248]={8'b00011000,
                 8'b00011000,
                 8'b00011000,
                 8'b00011000};
assign rom[249]={8'b00011000,
                 8'b00011000,
                 8'b00011000,
                 8'b00011000};

assign rom[250]={8'b00000000,
                 8'b01111110,
                 8'b01111000,
                 8'b01111100};
assign rom[251]={8'b01101110,
                 8'b01100110,
                 8'b00000110,
                 8'b00000000};

assign rom[252]={8'b00001000,
                 8'b00011000,
                 8'b00111000,
                 8'b01111000};
assign rom[253]={8'b00111000,
                 8'b00011000,
                 8'b00001000,
                 8'b00000000};

assign rom[254]={8'b00010000,
                 8'b00011000,
                 8'b00011100,
                 8'b00011110};
assign rom[255]={8'b00011100,
                 8'b00011000,
                 8'b00010000,
                 8'b00000000};
endmodule 
