


// Bit by Bit Multiply & Divide + Modulus
// Copyright © 2022 by Gregory Scott Callen
// All Rights Reserved.

// Migration from JavaScript to Verilog.

module mul (
   input wire        t,
   input wire [59:0] a,
   input wire [59:0] b,
   output reg [59:0] p
);

   // p = a * b

   p = 60'h0;

   always @ ( posedge t ) begin
      p = a [ 0 ] & b [ 0 ] ? p + ( 60'h1 << 0 ) : p ;
      p = a [ 0 ] & b [ 1 ] ? p + ( 60'h1 << 1 ) : p ;
      p = a [ 0 ] & b [ 2 ] ? p + ( 60'h1 << 2 ) : p ;
      p = a [ 0 ] & b [ 3 ] ? p + ( 60'h1 << 3 ) : p ;
      p = a [ 0 ] & b [ 4 ] ? p + ( 60'h1 << 4 ) : p ;
      p = a [ 0 ] & b [ 5 ] ? p + ( 60'h1 << 5 ) : p ;
      p = a [ 0 ] & b [ 6 ] ? p + ( 60'h1 << 6 ) : p ;
      p = a [ 0 ] & b [ 7 ] ? p + ( 60'h1 << 7 ) : p ;
      p = a [ 0 ] & b [ 8 ] ? p + ( 60'h1 << 8 ) : p ;
      p = a [ 0 ] & b [ 9 ] ? p + ( 60'h1 << 9 ) : p ;
      p = a [ 0 ] & b [ 10 ] ? p + ( 60'h1 << 10 ) : p ;
      p = a [ 0 ] & b [ 11 ] ? p + ( 60'h1 << 11 ) : p ;
      p = a [ 0 ] & b [ 12 ] ? p + ( 60'h1 << 12 ) : p ;
      p = a [ 0 ] & b [ 13 ] ? p + ( 60'h1 << 13 ) : p ;
      p = a [ 0 ] & b [ 14 ] ? p + ( 60'h1 << 14 ) : p ;
      p = a [ 0 ] & b [ 15 ] ? p + ( 60'h1 << 15 ) : p ;
      p = a [ 0 ] & b [ 16 ] ? p + ( 60'h1 << 16 ) : p ;
      p = a [ 0 ] & b [ 17 ] ? p + ( 60'h1 << 17 ) : p ;
      p = a [ 0 ] & b [ 18 ] ? p + ( 60'h1 << 18 ) : p ;
      p = a [ 0 ] & b [ 19 ] ? p + ( 60'h1 << 19 ) : p ;
      p = a [ 0 ] & b [ 20 ] ? p + ( 60'h1 << 20 ) : p ;
      p = a [ 0 ] & b [ 21 ] ? p + ( 60'h1 << 21 ) : p ;
      p = a [ 0 ] & b [ 22 ] ? p + ( 60'h1 << 22 ) : p ;
      p = a [ 0 ] & b [ 23 ] ? p + ( 60'h1 << 23 ) : p ;
      p = a [ 0 ] & b [ 24 ] ? p + ( 60'h1 << 24 ) : p ;
      p = a [ 0 ] & b [ 25 ] ? p + ( 60'h1 << 25 ) : p ;
      p = a [ 0 ] & b [ 26 ] ? p + ( 60'h1 << 26 ) : p ;
      p = a [ 0 ] & b [ 27 ] ? p + ( 60'h1 << 27 ) : p ;
      p = a [ 0 ] & b [ 28 ] ? p + ( 60'h1 << 28 ) : p ;
      p = a [ 0 ] & b [ 29 ] ? p + ( 60'h1 << 29 ) : p ;
      p = a [ 0 ] & b [ 30 ] ? p + ( 60'h1 << 30 ) : p ;
      p = a [ 0 ] & b [ 31 ] ? p + ( 60'h1 << 31 ) : p ;
      p = a [ 0 ] & b [ 32 ] ? p + ( 60'h1 << 32 ) : p ;
      p = a [ 0 ] & b [ 33 ] ? p + ( 60'h1 << 33 ) : p ;
      p = a [ 0 ] & b [ 34 ] ? p + ( 60'h1 << 34 ) : p ;
      p = a [ 0 ] & b [ 35 ] ? p + ( 60'h1 << 35 ) : p ;
      p = a [ 0 ] & b [ 36 ] ? p + ( 60'h1 << 36 ) : p ;
      p = a [ 0 ] & b [ 37 ] ? p + ( 60'h1 << 37 ) : p ;
      p = a [ 0 ] & b [ 38 ] ? p + ( 60'h1 << 38 ) : p ;
      p = a [ 0 ] & b [ 39 ] ? p + ( 60'h1 << 39 ) : p ;
      p = a [ 0 ] & b [ 40 ] ? p + ( 60'h1 << 40 ) : p ;
      p = a [ 0 ] & b [ 41 ] ? p + ( 60'h1 << 41 ) : p ;
      p = a [ 0 ] & b [ 42 ] ? p + ( 60'h1 << 42 ) : p ;
      p = a [ 0 ] & b [ 43 ] ? p + ( 60'h1 << 43 ) : p ;
      p = a [ 0 ] & b [ 44 ] ? p + ( 60'h1 << 44 ) : p ;
      p = a [ 0 ] & b [ 45 ] ? p + ( 60'h1 << 45 ) : p ;
      p = a [ 0 ] & b [ 46 ] ? p + ( 60'h1 << 46 ) : p ;
      p = a [ 0 ] & b [ 47 ] ? p + ( 60'h1 << 47 ) : p ;
      p = a [ 0 ] & b [ 48 ] ? p + ( 60'h1 << 48 ) : p ;
      p = a [ 0 ] & b [ 49 ] ? p + ( 60'h1 << 49 ) : p ;
      p = a [ 0 ] & b [ 50 ] ? p + ( 60'h1 << 50 ) : p ;
      p = a [ 0 ] & b [ 51 ] ? p + ( 60'h1 << 51 ) : p ;
      p = a [ 0 ] & b [ 52 ] ? p + ( 60'h1 << 52 ) : p ;
      p = a [ 0 ] & b [ 53 ] ? p + ( 60'h1 << 53 ) : p ;
      p = a [ 0 ] & b [ 54 ] ? p + ( 60'h1 << 54 ) : p ;
      p = a [ 0 ] & b [ 55 ] ? p + ( 60'h1 << 55 ) : p ;
      p = a [ 0 ] & b [ 56 ] ? p + ( 60'h1 << 56 ) : p ;
      p = a [ 0 ] & b [ 57 ] ? p + ( 60'h1 << 57 ) : p ;
      p = a [ 0 ] & b [ 58 ] ? p + ( 60'h1 << 58 ) : p ;
      p = a [ 0 ] & b [ 59 ] ? p + ( 60'h1 << 59 ) : p ;

// Bit by Bit Multiply & Divide + Modulus
// Copyright © 2022 by Gregory Scott Callen
// All Rights Reserved.

      p = a [ 1 ] & b [ 0 ] ? p + ( 60'h1 << 1 ) : p ;
      p = a [ 1 ] & b [ 1 ] ? p + ( 60'h1 << 2 ) : p ;
      p = a [ 1 ] & b [ 2 ] ? p + ( 60'h1 << 3 ) : p ;
      p = a [ 1 ] & b [ 3 ] ? p + ( 60'h1 << 4 ) : p ;
      p = a [ 1 ] & b [ 4 ] ? p + ( 60'h1 << 5 ) : p ;
      p = a [ 1 ] & b [ 5 ] ? p + ( 60'h1 << 6 ) : p ;
      p = a [ 1 ] & b [ 6 ] ? p + ( 60'h1 << 7 ) : p ;
      p = a [ 1 ] & b [ 7 ] ? p + ( 60'h1 << 8 ) : p ;
      p = a [ 1 ] & b [ 8 ] ? p + ( 60'h1 << 9 ) : p ;
      p = a [ 1 ] & b [ 9 ] ? p + ( 60'h1 << 10 ) : p ;
      p = a [ 1 ] & b [ 10 ] ? p + ( 60'h1 << 11 ) : p ;
      p = a [ 1 ] & b [ 11 ] ? p + ( 60'h1 << 12 ) : p ;
      p = a [ 1 ] & b [ 12 ] ? p + ( 60'h1 << 13 ) : p ;
      p = a [ 1 ] & b [ 13 ] ? p + ( 60'h1 << 14 ) : p ;
      p = a [ 1 ] & b [ 14 ] ? p + ( 60'h1 << 15 ) : p ;
      p = a [ 1 ] & b [ 15 ] ? p + ( 60'h1 << 16 ) : p ;
      p = a [ 1 ] & b [ 16 ] ? p + ( 60'h1 << 17 ) : p ;
      p = a [ 1 ] & b [ 17 ] ? p + ( 60'h1 << 18 ) : p ;
      p = a [ 1 ] & b [ 18 ] ? p + ( 60'h1 << 19 ) : p ;
      p = a [ 1 ] & b [ 19 ] ? p + ( 60'h1 << 20 ) : p ;
      p = a [ 1 ] & b [ 20 ] ? p + ( 60'h1 << 21 ) : p ;
      p = a [ 1 ] & b [ 21 ] ? p + ( 60'h1 << 22 ) : p ;
      p = a [ 1 ] & b [ 22 ] ? p + ( 60'h1 << 23 ) : p ;
      p = a [ 1 ] & b [ 23 ] ? p + ( 60'h1 << 24 ) : p ;
      p = a [ 1 ] & b [ 24 ] ? p + ( 60'h1 << 25 ) : p ;
      p = a [ 1 ] & b [ 25 ] ? p + ( 60'h1 << 26 ) : p ;
      p = a [ 1 ] & b [ 26 ] ? p + ( 60'h1 << 27 ) : p ;
      p = a [ 1 ] & b [ 27 ] ? p + ( 60'h1 << 28 ) : p ;
      p = a [ 1 ] & b [ 28 ] ? p + ( 60'h1 << 29 ) : p ;
      p = a [ 1 ] & b [ 29 ] ? p + ( 60'h1 << 30 ) : p ;
      p = a [ 1 ] & b [ 30 ] ? p + ( 60'h1 << 31 ) : p ;
      p = a [ 1 ] & b [ 31 ] ? p + ( 60'h1 << 32 ) : p ;
      p = a [ 1 ] & b [ 32 ] ? p + ( 60'h1 << 33 ) : p ;
      p = a [ 1 ] & b [ 33 ] ? p + ( 60'h1 << 34 ) : p ;
      p = a [ 1 ] & b [ 34 ] ? p + ( 60'h1 << 35 ) : p ;
      p = a [ 1 ] & b [ 35 ] ? p + ( 60'h1 << 36 ) : p ;
      p = a [ 1 ] & b [ 36 ] ? p + ( 60'h1 << 37 ) : p ;
      p = a [ 1 ] & b [ 37 ] ? p + ( 60'h1 << 38 ) : p ;
      p = a [ 1 ] & b [ 38 ] ? p + ( 60'h1 << 39 ) : p ;
      p = a [ 1 ] & b [ 39 ] ? p + ( 60'h1 << 40 ) : p ;
      p = a [ 1 ] & b [ 40 ] ? p + ( 60'h1 << 41 ) : p ;
      p = a [ 1 ] & b [ 41 ] ? p + ( 60'h1 << 42 ) : p ;
      p = a [ 1 ] & b [ 42 ] ? p + ( 60'h1 << 43 ) : p ;
      p = a [ 1 ] & b [ 43 ] ? p + ( 60'h1 << 44 ) : p ;
      p = a [ 1 ] & b [ 44 ] ? p + ( 60'h1 << 45 ) : p ;
      p = a [ 1 ] & b [ 45 ] ? p + ( 60'h1 << 46 ) : p ;
      p = a [ 1 ] & b [ 46 ] ? p + ( 60'h1 << 47 ) : p ;
      p = a [ 1 ] & b [ 47 ] ? p + ( 60'h1 << 48 ) : p ;
      p = a [ 1 ] & b [ 48 ] ? p + ( 60'h1 << 49 ) : p ;
      p = a [ 1 ] & b [ 49 ] ? p + ( 60'h1 << 50 ) : p ;
      p = a [ 1 ] & b [ 50 ] ? p + ( 60'h1 << 51 ) : p ;
      p = a [ 1 ] & b [ 51 ] ? p + ( 60'h1 << 52 ) : p ;
      p = a [ 1 ] & b [ 52 ] ? p + ( 60'h1 << 53 ) : p ;
      p = a [ 1 ] & b [ 53 ] ? p + ( 60'h1 << 54 ) : p ;
      p = a [ 1 ] & b [ 54 ] ? p + ( 60'h1 << 55 ) : p ;
      p = a [ 1 ] & b [ 55 ] ? p + ( 60'h1 << 56 ) : p ;
      p = a [ 1 ] & b [ 56 ] ? p + ( 60'h1 << 57 ) : p ;
      p = a [ 1 ] & b [ 57 ] ? p + ( 60'h1 << 58 ) : p ;
      p = a [ 1 ] & b [ 58 ] ? p + ( 60'h1 << 59 ) : p ;

// Bit by Bit Multiply & Divide + Modulus
// Copyright © 2022 by Gregory Scott Callen
// All Rights Reserved.

      p = a [ 2 ] & b [ 0 ] ? p + ( 60'h1 << 2 ) : p ;
      p = a [ 2 ] & b [ 1 ] ? p + ( 60'h1 << 3 ) : p ;
      p = a [ 2 ] & b [ 2 ] ? p + ( 60'h1 << 4 ) : p ;
      p = a [ 2 ] & b [ 3 ] ? p + ( 60'h1 << 5 ) : p ;
      p = a [ 2 ] & b [ 4 ] ? p + ( 60'h1 << 6 ) : p ;
      p = a [ 2 ] & b [ 5 ] ? p + ( 60'h1 << 7 ) : p ;
      p = a [ 2 ] & b [ 6 ] ? p + ( 60'h1 << 8 ) : p ;
      p = a [ 2 ] & b [ 7 ] ? p + ( 60'h1 << 9 ) : p ;
      p = a [ 2 ] & b [ 8 ] ? p + ( 60'h1 << 10 ) : p ;
      p = a [ 2 ] & b [ 9 ] ? p + ( 60'h1 << 11 ) : p ;
      p = a [ 2 ] & b [ 10 ] ? p + ( 60'h1 << 12 ) : p ;
      p = a [ 2 ] & b [ 11 ] ? p + ( 60'h1 << 13 ) : p ;
      p = a [ 2 ] & b [ 12 ] ? p + ( 60'h1 << 14 ) : p ;
      p = a [ 2 ] & b [ 13 ] ? p + ( 60'h1 << 15 ) : p ;
      p = a [ 2 ] & b [ 14 ] ? p + ( 60'h1 << 16 ) : p ;
      p = a [ 2 ] & b [ 15 ] ? p + ( 60'h1 << 17 ) : p ;
      p = a [ 2 ] & b [ 16 ] ? p + ( 60'h1 << 18 ) : p ;
      p = a [ 2 ] & b [ 17 ] ? p + ( 60'h1 << 19 ) : p ;
      p = a [ 2 ] & b [ 18 ] ? p + ( 60'h1 << 20 ) : p ;
      p = a [ 2 ] & b [ 19 ] ? p + ( 60'h1 << 21 ) : p ;
      p = a [ 2 ] & b [ 20 ] ? p + ( 60'h1 << 22 ) : p ;
      p = a [ 2 ] & b [ 21 ] ? p + ( 60'h1 << 23 ) : p ;
      p = a [ 2 ] & b [ 22 ] ? p + ( 60'h1 << 24 ) : p ;
      p = a [ 2 ] & b [ 23 ] ? p + ( 60'h1 << 25 ) : p ;
      p = a [ 2 ] & b [ 24 ] ? p + ( 60'h1 << 26 ) : p ;
      p = a [ 2 ] & b [ 25 ] ? p + ( 60'h1 << 27 ) : p ;
      p = a [ 2 ] & b [ 26 ] ? p + ( 60'h1 << 28 ) : p ;
      p = a [ 2 ] & b [ 27 ] ? p + ( 60'h1 << 29 ) : p ;
      p = a [ 2 ] & b [ 28 ] ? p + ( 60'h1 << 30 ) : p ;
      p = a [ 2 ] & b [ 29 ] ? p + ( 60'h1 << 31 ) : p ;
      p = a [ 2 ] & b [ 30 ] ? p + ( 60'h1 << 32 ) : p ;
      p = a [ 2 ] & b [ 31 ] ? p + ( 60'h1 << 33 ) : p ;
      p = a [ 2 ] & b [ 32 ] ? p + ( 60'h1 << 34 ) : p ;
      p = a [ 2 ] & b [ 33 ] ? p + ( 60'h1 << 35 ) : p ;
      p = a [ 2 ] & b [ 34 ] ? p + ( 60'h1 << 36 ) : p ;
      p = a [ 2 ] & b [ 35 ] ? p + ( 60'h1 << 37 ) : p ;
      p = a [ 2 ] & b [ 36 ] ? p + ( 60'h1 << 38 ) : p ;
      p = a [ 2 ] & b [ 37 ] ? p + ( 60'h1 << 39 ) : p ;
      p = a [ 2 ] & b [ 38 ] ? p + ( 60'h1 << 40 ) : p ;
      p = a [ 2 ] & b [ 39 ] ? p + ( 60'h1 << 41 ) : p ;
      p = a [ 2 ] & b [ 40 ] ? p + ( 60'h1 << 42 ) : p ;
      p = a [ 2 ] & b [ 41 ] ? p + ( 60'h1 << 43 ) : p ;
      p = a [ 2 ] & b [ 42 ] ? p + ( 60'h1 << 44 ) : p ;
      p = a [ 2 ] & b [ 43 ] ? p + ( 60'h1 << 45 ) : p ;
      p = a [ 2 ] & b [ 44 ] ? p + ( 60'h1 << 46 ) : p ;
      p = a [ 2 ] & b [ 45 ] ? p + ( 60'h1 << 47 ) : p ;
      p = a [ 2 ] & b [ 46 ] ? p + ( 60'h1 << 48 ) : p ;
      p = a [ 2 ] & b [ 47 ] ? p + ( 60'h1 << 49 ) : p ;
      p = a [ 2 ] & b [ 48 ] ? p + ( 60'h1 << 50 ) : p ;
      p = a [ 2 ] & b [ 49 ] ? p + ( 60'h1 << 51 ) : p ;
      p = a [ 2 ] & b [ 50 ] ? p + ( 60'h1 << 52 ) : p ;
      p = a [ 2 ] & b [ 51 ] ? p + ( 60'h1 << 53 ) : p ;
      p = a [ 2 ] & b [ 52 ] ? p + ( 60'h1 << 54 ) : p ;
      p = a [ 2 ] & b [ 53 ] ? p + ( 60'h1 << 55 ) : p ;
      p = a [ 2 ] & b [ 54 ] ? p + ( 60'h1 << 56 ) : p ;
      p = a [ 2 ] & b [ 55 ] ? p + ( 60'h1 << 57 ) : p ;
      p = a [ 2 ] & b [ 56 ] ? p + ( 60'h1 << 58 ) : p ;
      p = a [ 2 ] & b [ 57 ] ? p + ( 60'h1 << 59 ) : p ;

// Bit by Bit Multiply & Divide + Modulus
// Copyright © 2022 by Gregory Scott Callen
// All Rights Reserved.

      p = a [ 3 ] & b [ 0 ] ? p + ( 60'h1 << 3 ) : p ;
      p = a [ 3 ] & b [ 1 ] ? p + ( 60'h1 << 4 ) : p ;
      p = a [ 3 ] & b [ 2 ] ? p + ( 60'h1 << 5 ) : p ;
      p = a [ 3 ] & b [ 3 ] ? p + ( 60'h1 << 6 ) : p ;
      p = a [ 3 ] & b [ 4 ] ? p + ( 60'h1 << 7 ) : p ;
      p = a [ 3 ] & b [ 5 ] ? p + ( 60'h1 << 8 ) : p ;
      p = a [ 3 ] & b [ 6 ] ? p + ( 60'h1 << 9 ) : p ;
      p = a [ 3 ] & b [ 7 ] ? p + ( 60'h1 << 10 ) : p ;
      p = a [ 3 ] & b [ 8 ] ? p + ( 60'h1 << 11 ) : p ;
      p = a [ 3 ] & b [ 9 ] ? p + ( 60'h1 << 12 ) : p ;
      p = a [ 3 ] & b [ 10 ] ? p + ( 60'h1 << 13 ) : p ;
      p = a [ 3 ] & b [ 11 ] ? p + ( 60'h1 << 14 ) : p ;
      p = a [ 3 ] & b [ 12 ] ? p + ( 60'h1 << 15 ) : p ;
      p = a [ 3 ] & b [ 13 ] ? p + ( 60'h1 << 16 ) : p ;
      p = a [ 3 ] & b [ 14 ] ? p + ( 60'h1 << 17 ) : p ;
      p = a [ 3 ] & b [ 15 ] ? p + ( 60'h1 << 18 ) : p ;
      p = a [ 3 ] & b [ 16 ] ? p + ( 60'h1 << 19 ) : p ;
      p = a [ 3 ] & b [ 17 ] ? p + ( 60'h1 << 20 ) : p ;
      p = a [ 3 ] & b [ 18 ] ? p + ( 60'h1 << 21 ) : p ;
      p = a [ 3 ] & b [ 19 ] ? p + ( 60'h1 << 22 ) : p ;
      p = a [ 3 ] & b [ 20 ] ? p + ( 60'h1 << 23 ) : p ;
      p = a [ 3 ] & b [ 21 ] ? p + ( 60'h1 << 24 ) : p ;
      p = a [ 3 ] & b [ 22 ] ? p + ( 60'h1 << 25 ) : p ;
      p = a [ 3 ] & b [ 23 ] ? p + ( 60'h1 << 26 ) : p ;
      p = a [ 3 ] & b [ 24 ] ? p + ( 60'h1 << 27 ) : p ;
      p = a [ 3 ] & b [ 25 ] ? p + ( 60'h1 << 28 ) : p ;
      p = a [ 3 ] & b [ 26 ] ? p + ( 60'h1 << 29 ) : p ;
      p = a [ 3 ] & b [ 27 ] ? p + ( 60'h1 << 30 ) : p ;
      p = a [ 3 ] & b [ 28 ] ? p + ( 60'h1 << 31 ) : p ;
      p = a [ 3 ] & b [ 29 ] ? p + ( 60'h1 << 32 ) : p ;
      p = a [ 3 ] & b [ 30 ] ? p + ( 60'h1 << 33 ) : p ;
      p = a [ 3 ] & b [ 31 ] ? p + ( 60'h1 << 34 ) : p ;
      p = a [ 3 ] & b [ 32 ] ? p + ( 60'h1 << 35 ) : p ;
      p = a [ 3 ] & b [ 33 ] ? p + ( 60'h1 << 36 ) : p ;
      p = a [ 3 ] & b [ 34 ] ? p + ( 60'h1 << 37 ) : p ;
      p = a [ 3 ] & b [ 35 ] ? p + ( 60'h1 << 38 ) : p ;
      p = a [ 3 ] & b [ 36 ] ? p + ( 60'h1 << 39 ) : p ;
      p = a [ 3 ] & b [ 37 ] ? p + ( 60'h1 << 40 ) : p ;
      p = a [ 3 ] & b [ 38 ] ? p + ( 60'h1 << 41 ) : p ;
      p = a [ 3 ] & b [ 39 ] ? p + ( 60'h1 << 42 ) : p ;
      p = a [ 3 ] & b [ 40 ] ? p + ( 60'h1 << 43 ) : p ;
      p = a [ 3 ] & b [ 41 ] ? p + ( 60'h1 << 44 ) : p ;
      p = a [ 3 ] & b [ 42 ] ? p + ( 60'h1 << 45 ) : p ;
      p = a [ 3 ] & b [ 43 ] ? p + ( 60'h1 << 46 ) : p ;
      p = a [ 3 ] & b [ 44 ] ? p + ( 60'h1 << 47 ) : p ;
      p = a [ 3 ] & b [ 45 ] ? p + ( 60'h1 << 48 ) : p ;
      p = a [ 3 ] & b [ 46 ] ? p + ( 60'h1 << 49 ) : p ;
      p = a [ 3 ] & b [ 47 ] ? p + ( 60'h1 << 50 ) : p ;
      p = a [ 3 ] & b [ 48 ] ? p + ( 60'h1 << 51 ) : p ;
      p = a [ 3 ] & b [ 49 ] ? p + ( 60'h1 << 52 ) : p ;
      p = a [ 3 ] & b [ 50 ] ? p + ( 60'h1 << 53 ) : p ;
      p = a [ 3 ] & b [ 51 ] ? p + ( 60'h1 << 54 ) : p ;
      p = a [ 3 ] & b [ 52 ] ? p + ( 60'h1 << 55 ) : p ;
      p = a [ 3 ] & b [ 53 ] ? p + ( 60'h1 << 56 ) : p ;
      p = a [ 3 ] & b [ 54 ] ? p + ( 60'h1 << 57 ) : p ;
      p = a [ 3 ] & b [ 55 ] ? p + ( 60'h1 << 58 ) : p ;
      p = a [ 3 ] & b [ 56 ] ? p + ( 60'h1 << 59 ) : p ;

// Bit by Bit Multiply & Divide + Modulus
// Copyright © 2022 by Gregory Scott Callen
// All Rights Reserved.

      p = a [ 4 ] & b [ 0 ] ? p + ( 60'h1 << 4 ) : p ;
      p = a [ 4 ] & b [ 1 ] ? p + ( 60'h1 << 5 ) : p ;
      p = a [ 4 ] & b [ 2 ] ? p + ( 60'h1 << 6 ) : p ;
      p = a [ 4 ] & b [ 3 ] ? p + ( 60'h1 << 7 ) : p ;
      p = a [ 4 ] & b [ 4 ] ? p + ( 60'h1 << 8 ) : p ;
      p = a [ 4 ] & b [ 5 ] ? p + ( 60'h1 << 9 ) : p ;
      p = a [ 4 ] & b [ 6 ] ? p + ( 60'h1 << 10 ) : p ;
      p = a [ 4 ] & b [ 7 ] ? p + ( 60'h1 << 11 ) : p ;
      p = a [ 4 ] & b [ 8 ] ? p + ( 60'h1 << 12 ) : p ;
      p = a [ 4 ] & b [ 9 ] ? p + ( 60'h1 << 13 ) : p ;
      p = a [ 4 ] & b [ 10 ] ? p + ( 60'h1 << 14 ) : p ;
      p = a [ 4 ] & b [ 11 ] ? p + ( 60'h1 << 15 ) : p ;
      p = a [ 4 ] & b [ 12 ] ? p + ( 60'h1 << 16 ) : p ;
      p = a [ 4 ] & b [ 13 ] ? p + ( 60'h1 << 17 ) : p ;
      p = a [ 4 ] & b [ 14 ] ? p + ( 60'h1 << 18 ) : p ;
      p = a [ 4 ] & b [ 15 ] ? p + ( 60'h1 << 19 ) : p ;
      p = a [ 4 ] & b [ 16 ] ? p + ( 60'h1 << 20 ) : p ;
      p = a [ 4 ] & b [ 17 ] ? p + ( 60'h1 << 21 ) : p ;
      p = a [ 4 ] & b [ 18 ] ? p + ( 60'h1 << 22 ) : p ;
      p = a [ 4 ] & b [ 19 ] ? p + ( 60'h1 << 23 ) : p ;
      p = a [ 4 ] & b [ 20 ] ? p + ( 60'h1 << 24 ) : p ;
      p = a [ 4 ] & b [ 21 ] ? p + ( 60'h1 << 25 ) : p ;
      p = a [ 4 ] & b [ 22 ] ? p + ( 60'h1 << 26 ) : p ;
      p = a [ 4 ] & b [ 23 ] ? p + ( 60'h1 << 27 ) : p ;
      p = a [ 4 ] & b [ 24 ] ? p + ( 60'h1 << 28 ) : p ;
      p = a [ 4 ] & b [ 25 ] ? p + ( 60'h1 << 29 ) : p ;
      p = a [ 4 ] & b [ 26 ] ? p + ( 60'h1 << 30 ) : p ;
      p = a [ 4 ] & b [ 27 ] ? p + ( 60'h1 << 31 ) : p ;
      p = a [ 4 ] & b [ 28 ] ? p + ( 60'h1 << 32 ) : p ;
      p = a [ 4 ] & b [ 29 ] ? p + ( 60'h1 << 33 ) : p ;
      p = a [ 4 ] & b [ 30 ] ? p + ( 60'h1 << 34 ) : p ;
      p = a [ 4 ] & b [ 31 ] ? p + ( 60'h1 << 35 ) : p ;
      p = a [ 4 ] & b [ 32 ] ? p + ( 60'h1 << 36 ) : p ;
      p = a [ 4 ] & b [ 33 ] ? p + ( 60'h1 << 37 ) : p ;
      p = a [ 4 ] & b [ 34 ] ? p + ( 60'h1 << 38 ) : p ;
      p = a [ 4 ] & b [ 35 ] ? p + ( 60'h1 << 39 ) : p ;
      p = a [ 4 ] & b [ 36 ] ? p + ( 60'h1 << 40 ) : p ;
      p = a [ 4 ] & b [ 37 ] ? p + ( 60'h1 << 41 ) : p ;
      p = a [ 4 ] & b [ 38 ] ? p + ( 60'h1 << 42 ) : p ;
      p = a [ 4 ] & b [ 39 ] ? p + ( 60'h1 << 43 ) : p ;
      p = a [ 4 ] & b [ 40 ] ? p + ( 60'h1 << 44 ) : p ;
      p = a [ 4 ] & b [ 41 ] ? p + ( 60'h1 << 45 ) : p ;
      p = a [ 4 ] & b [ 42 ] ? p + ( 60'h1 << 46 ) : p ;
      p = a [ 4 ] & b [ 43 ] ? p + ( 60'h1 << 47 ) : p ;
      p = a [ 4 ] & b [ 44 ] ? p + ( 60'h1 << 48 ) : p ;
      p = a [ 4 ] & b [ 45 ] ? p + ( 60'h1 << 49 ) : p ;
      p = a [ 4 ] & b [ 46 ] ? p + ( 60'h1 << 50 ) : p ;
      p = a [ 4 ] & b [ 47 ] ? p + ( 60'h1 << 51 ) : p ;
      p = a [ 4 ] & b [ 48 ] ? p + ( 60'h1 << 52 ) : p ;
      p = a [ 4 ] & b [ 49 ] ? p + ( 60'h1 << 53 ) : p ;
      p = a [ 4 ] & b [ 50 ] ? p + ( 60'h1 << 54 ) : p ;
      p = a [ 4 ] & b [ 51 ] ? p + ( 60'h1 << 55 ) : p ;
      p = a [ 4 ] & b [ 52 ] ? p + ( 60'h1 << 56 ) : p ;
      p = a [ 4 ] & b [ 53 ] ? p + ( 60'h1 << 57 ) : p ;
      p = a [ 4 ] & b [ 54 ] ? p + ( 60'h1 << 58 ) : p ;
      p = a [ 4 ] & b [ 55 ] ? p + ( 60'h1 << 59 ) : p ;

// Bit by Bit Multiply & Divide + Modulus
// Copyright © 2022 by Gregory Scott Callen
// All Rights Reserved.

      p = a [ 5 ] & b [ 0 ] ? p + ( 60'h1 << 5 ) : p ;
      p = a [ 5 ] & b [ 1 ] ? p + ( 60'h1 << 6 ) : p ;
      p = a [ 5 ] & b [ 2 ] ? p + ( 60'h1 << 7 ) : p ;
      p = a [ 5 ] & b [ 3 ] ? p + ( 60'h1 << 8 ) : p ;
      p = a [ 5 ] & b [ 4 ] ? p + ( 60'h1 << 9 ) : p ;
      p = a [ 5 ] & b [ 5 ] ? p + ( 60'h1 << 10 ) : p ;
      p = a [ 5 ] & b [ 6 ] ? p + ( 60'h1 << 11 ) : p ;
      p = a [ 5 ] & b [ 7 ] ? p + ( 60'h1 << 12 ) : p ;
      p = a [ 5 ] & b [ 8 ] ? p + ( 60'h1 << 13 ) : p ;
      p = a [ 5 ] & b [ 9 ] ? p + ( 60'h1 << 14 ) : p ;
      p = a [ 5 ] & b [ 10 ] ? p + ( 60'h1 << 15 ) : p ;
      p = a [ 5 ] & b [ 11 ] ? p + ( 60'h1 << 16 ) : p ;
      p = a [ 5 ] & b [ 12 ] ? p + ( 60'h1 << 17 ) : p ;
      p = a [ 5 ] & b [ 13 ] ? p + ( 60'h1 << 18 ) : p ;
      p = a [ 5 ] & b [ 14 ] ? p + ( 60'h1 << 19 ) : p ;
      p = a [ 5 ] & b [ 15 ] ? p + ( 60'h1 << 20 ) : p ;
      p = a [ 5 ] & b [ 16 ] ? p + ( 60'h1 << 21 ) : p ;
      p = a [ 5 ] & b [ 17 ] ? p + ( 60'h1 << 22 ) : p ;
      p = a [ 5 ] & b [ 18 ] ? p + ( 60'h1 << 23 ) : p ;
      p = a [ 5 ] & b [ 19 ] ? p + ( 60'h1 << 24 ) : p ;
      p = a [ 5 ] & b [ 20 ] ? p + ( 60'h1 << 25 ) : p ;
      p = a [ 5 ] & b [ 21 ] ? p + ( 60'h1 << 26 ) : p ;
      p = a [ 5 ] & b [ 22 ] ? p + ( 60'h1 << 27 ) : p ;
      p = a [ 5 ] & b [ 23 ] ? p + ( 60'h1 << 28 ) : p ;
      p = a [ 5 ] & b [ 24 ] ? p + ( 60'h1 << 29 ) : p ;
      p = a [ 5 ] & b [ 25 ] ? p + ( 60'h1 << 30 ) : p ;
      p = a [ 5 ] & b [ 26 ] ? p + ( 60'h1 << 31 ) : p ;
      p = a [ 5 ] & b [ 27 ] ? p + ( 60'h1 << 32 ) : p ;
      p = a [ 5 ] & b [ 28 ] ? p + ( 60'h1 << 33 ) : p ;
      p = a [ 5 ] & b [ 29 ] ? p + ( 60'h1 << 34 ) : p ;
      p = a [ 5 ] & b [ 30 ] ? p + ( 60'h1 << 35 ) : p ;
      p = a [ 5 ] & b [ 31 ] ? p + ( 60'h1 << 36 ) : p ;
      p = a [ 5 ] & b [ 32 ] ? p + ( 60'h1 << 37 ) : p ;
      p = a [ 5 ] & b [ 33 ] ? p + ( 60'h1 << 38 ) : p ;
      p = a [ 5 ] & b [ 34 ] ? p + ( 60'h1 << 39 ) : p ;
      p = a [ 5 ] & b [ 35 ] ? p + ( 60'h1 << 40 ) : p ;
      p = a [ 5 ] & b [ 36 ] ? p + ( 60'h1 << 41 ) : p ;
      p = a [ 5 ] & b [ 37 ] ? p + ( 60'h1 << 42 ) : p ;
      p = a [ 5 ] & b [ 38 ] ? p + ( 60'h1 << 43 ) : p ;
      p = a [ 5 ] & b [ 39 ] ? p + ( 60'h1 << 44 ) : p ;
      p = a [ 5 ] & b [ 40 ] ? p + ( 60'h1 << 45 ) : p ;
      p = a [ 5 ] & b [ 41 ] ? p + ( 60'h1 << 46 ) : p ;
      p = a [ 5 ] & b [ 42 ] ? p + ( 60'h1 << 47 ) : p ;
      p = a [ 5 ] & b [ 43 ] ? p + ( 60'h1 << 48 ) : p ;
      p = a [ 5 ] & b [ 44 ] ? p + ( 60'h1 << 49 ) : p ;
      p = a [ 5 ] & b [ 45 ] ? p + ( 60'h1 << 50 ) : p ;
      p = a [ 5 ] & b [ 46 ] ? p + ( 60'h1 << 51 ) : p ;
      p = a [ 5 ] & b [ 47 ] ? p + ( 60'h1 << 52 ) : p ;
      p = a [ 5 ] & b [ 48 ] ? p + ( 60'h1 << 53 ) : p ;
      p = a [ 5 ] & b [ 49 ] ? p + ( 60'h1 << 54 ) : p ;
      p = a [ 5 ] & b [ 50 ] ? p + ( 60'h1 << 55 ) : p ;
      p = a [ 5 ] & b [ 51 ] ? p + ( 60'h1 << 56 ) : p ;
      p = a [ 5 ] & b [ 52 ] ? p + ( 60'h1 << 57 ) : p ;
      p = a [ 5 ] & b [ 53 ] ? p + ( 60'h1 << 58 ) : p ;
      p = a [ 5 ] & b [ 54 ] ? p + ( 60'h1 << 59 ) : p ;

// Bit by Bit Multiply & Divide + Modulus
// Copyright © 2022 by Gregory Scott Callen
// All Rights Reserved.

      p = a [ 6 ] & b [ 0 ] ? p + ( 60'h1 << 6 ) : p ;
      p = a [ 6 ] & b [ 1 ] ? p + ( 60'h1 << 7 ) : p ;
      p = a [ 6 ] & b [ 2 ] ? p + ( 60'h1 << 8 ) : p ;
      p = a [ 6 ] & b [ 3 ] ? p + ( 60'h1 << 9 ) : p ;
      p = a [ 6 ] & b [ 4 ] ? p + ( 60'h1 << 10 ) : p ;
      p = a [ 6 ] & b [ 5 ] ? p + ( 60'h1 << 11 ) : p ;
      p = a [ 6 ] & b [ 6 ] ? p + ( 60'h1 << 12 ) : p ;
      p = a [ 6 ] & b [ 7 ] ? p + ( 60'h1 << 13 ) : p ;
      p = a [ 6 ] & b [ 8 ] ? p + ( 60'h1 << 14 ) : p ;
      p = a [ 6 ] & b [ 9 ] ? p + ( 60'h1 << 15 ) : p ;
      p = a [ 6 ] & b [ 10 ] ? p + ( 60'h1 << 16 ) : p ;
      p = a [ 6 ] & b [ 11 ] ? p + ( 60'h1 << 17 ) : p ;
      p = a [ 6 ] & b [ 12 ] ? p + ( 60'h1 << 18 ) : p ;
      p = a [ 6 ] & b [ 13 ] ? p + ( 60'h1 << 19 ) : p ;
      p = a [ 6 ] & b [ 14 ] ? p + ( 60'h1 << 20 ) : p ;
      p = a [ 6 ] & b [ 15 ] ? p + ( 60'h1 << 21 ) : p ;
      p = a [ 6 ] & b [ 16 ] ? p + ( 60'h1 << 22 ) : p ;
      p = a [ 6 ] & b [ 17 ] ? p + ( 60'h1 << 23 ) : p ;
      p = a [ 6 ] & b [ 18 ] ? p + ( 60'h1 << 24 ) : p ;
      p = a [ 6 ] & b [ 19 ] ? p + ( 60'h1 << 25 ) : p ;
      p = a [ 6 ] & b [ 20 ] ? p + ( 60'h1 << 26 ) : p ;
      p = a [ 6 ] & b [ 21 ] ? p + ( 60'h1 << 27 ) : p ;
      p = a [ 6 ] & b [ 22 ] ? p + ( 60'h1 << 28 ) : p ;
      p = a [ 6 ] & b [ 23 ] ? p + ( 60'h1 << 29 ) : p ;
      p = a [ 6 ] & b [ 24 ] ? p + ( 60'h1 << 30 ) : p ;
      p = a [ 6 ] & b [ 25 ] ? p + ( 60'h1 << 31 ) : p ;
      p = a [ 6 ] & b [ 26 ] ? p + ( 60'h1 << 32 ) : p ;
      p = a [ 6 ] & b [ 27 ] ? p + ( 60'h1 << 33 ) : p ;
      p = a [ 6 ] & b [ 28 ] ? p + ( 60'h1 << 34 ) : p ;
      p = a [ 6 ] & b [ 29 ] ? p + ( 60'h1 << 35 ) : p ;
      p = a [ 6 ] & b [ 30 ] ? p + ( 60'h1 << 36 ) : p ;
      p = a [ 6 ] & b [ 31 ] ? p + ( 60'h1 << 37 ) : p ;
      p = a [ 6 ] & b [ 32 ] ? p + ( 60'h1 << 38 ) : p ;
      p = a [ 6 ] & b [ 33 ] ? p + ( 60'h1 << 39 ) : p ;
      p = a [ 6 ] & b [ 34 ] ? p + ( 60'h1 << 40 ) : p ;
      p = a [ 6 ] & b [ 35 ] ? p + ( 60'h1 << 41 ) : p ;
      p = a [ 6 ] & b [ 36 ] ? p + ( 60'h1 << 42 ) : p ;
      p = a [ 6 ] & b [ 37 ] ? p + ( 60'h1 << 43 ) : p ;
      p = a [ 6 ] & b [ 38 ] ? p + ( 60'h1 << 44 ) : p ;
      p = a [ 6 ] & b [ 39 ] ? p + ( 60'h1 << 45 ) : p ;
      p = a [ 6 ] & b [ 40 ] ? p + ( 60'h1 << 46 ) : p ;
      p = a [ 6 ] & b [ 41 ] ? p + ( 60'h1 << 47 ) : p ;
      p = a [ 6 ] & b [ 42 ] ? p + ( 60'h1 << 48 ) : p ;
      p = a [ 6 ] & b [ 43 ] ? p + ( 60'h1 << 49 ) : p ;
      p = a [ 6 ] & b [ 44 ] ? p + ( 60'h1 << 50 ) : p ;
      p = a [ 6 ] & b [ 45 ] ? p + ( 60'h1 << 51 ) : p ;
      p = a [ 6 ] & b [ 46 ] ? p + ( 60'h1 << 52 ) : p ;
      p = a [ 6 ] & b [ 47 ] ? p + ( 60'h1 << 53 ) : p ;
      p = a [ 6 ] & b [ 48 ] ? p + ( 60'h1 << 54 ) : p ;
      p = a [ 6 ] & b [ 49 ] ? p + ( 60'h1 << 55 ) : p ;
      p = a [ 6 ] & b [ 50 ] ? p + ( 60'h1 << 56 ) : p ;
      p = a [ 6 ] & b [ 51 ] ? p + ( 60'h1 << 57 ) : p ;
      p = a [ 6 ] & b [ 52 ] ? p + ( 60'h1 << 58 ) : p ;
      p = a [ 6 ] & b [ 53 ] ? p + ( 60'h1 << 59 ) : p ;

// Bit by Bit Multiply & Divide + Modulus
// Copyright © 2022 by Gregory Scott Callen
// All Rights Reserved.

      p = a [ 7 ] & b [ 0 ] ? p + ( 60'h1 << 7 ) : p ;
      p = a [ 7 ] & b [ 1 ] ? p + ( 60'h1 << 8 ) : p ;
      p = a [ 7 ] & b [ 2 ] ? p + ( 60'h1 << 9 ) : p ;
      p = a [ 7 ] & b [ 3 ] ? p + ( 60'h1 << 10 ) : p ;
      p = a [ 7 ] & b [ 4 ] ? p + ( 60'h1 << 11 ) : p ;
      p = a [ 7 ] & b [ 5 ] ? p + ( 60'h1 << 12 ) : p ;
      p = a [ 7 ] & b [ 6 ] ? p + ( 60'h1 << 13 ) : p ;
      p = a [ 7 ] & b [ 7 ] ? p + ( 60'h1 << 14 ) : p ;
      p = a [ 7 ] & b [ 8 ] ? p + ( 60'h1 << 15 ) : p ;
      p = a [ 7 ] & b [ 9 ] ? p + ( 60'h1 << 16 ) : p ;
      p = a [ 7 ] & b [ 10 ] ? p + ( 60'h1 << 17 ) : p ;
      p = a [ 7 ] & b [ 11 ] ? p + ( 60'h1 << 18 ) : p ;
      p = a [ 7 ] & b [ 12 ] ? p + ( 60'h1 << 19 ) : p ;
      p = a [ 7 ] & b [ 13 ] ? p + ( 60'h1 << 20 ) : p ;
      p = a [ 7 ] & b [ 14 ] ? p + ( 60'h1 << 21 ) : p ;
      p = a [ 7 ] & b [ 15 ] ? p + ( 60'h1 << 22 ) : p ;
      p = a [ 7 ] & b [ 16 ] ? p + ( 60'h1 << 23 ) : p ;
      p = a [ 7 ] & b [ 17 ] ? p + ( 60'h1 << 24 ) : p ;
      p = a [ 7 ] & b [ 18 ] ? p + ( 60'h1 << 25 ) : p ;
      p = a [ 7 ] & b [ 19 ] ? p + ( 60'h1 << 26 ) : p ;
      p = a [ 7 ] & b [ 20 ] ? p + ( 60'h1 << 27 ) : p ;
      p = a [ 7 ] & b [ 21 ] ? p + ( 60'h1 << 28 ) : p ;
      p = a [ 7 ] & b [ 22 ] ? p + ( 60'h1 << 29 ) : p ;
      p = a [ 7 ] & b [ 23 ] ? p + ( 60'h1 << 30 ) : p ;
      p = a [ 7 ] & b [ 24 ] ? p + ( 60'h1 << 31 ) : p ;
      p = a [ 7 ] & b [ 25 ] ? p + ( 60'h1 << 32 ) : p ;
      p = a [ 7 ] & b [ 26 ] ? p + ( 60'h1 << 33 ) : p ;
      p = a [ 7 ] & b [ 27 ] ? p + ( 60'h1 << 34 ) : p ;
      p = a [ 7 ] & b [ 28 ] ? p + ( 60'h1 << 35 ) : p ;
      p = a [ 7 ] & b [ 29 ] ? p + ( 60'h1 << 36 ) : p ;
      p = a [ 7 ] & b [ 30 ] ? p + ( 60'h1 << 37 ) : p ;
      p = a [ 7 ] & b [ 31 ] ? p + ( 60'h1 << 38 ) : p ;
      p = a [ 7 ] & b [ 32 ] ? p + ( 60'h1 << 39 ) : p ;
      p = a [ 7 ] & b [ 33 ] ? p + ( 60'h1 << 40 ) : p ;
      p = a [ 7 ] & b [ 34 ] ? p + ( 60'h1 << 41 ) : p ;
      p = a [ 7 ] & b [ 35 ] ? p + ( 60'h1 << 42 ) : p ;
      p = a [ 7 ] & b [ 36 ] ? p + ( 60'h1 << 43 ) : p ;
      p = a [ 7 ] & b [ 37 ] ? p + ( 60'h1 << 44 ) : p ;
      p = a [ 7 ] & b [ 38 ] ? p + ( 60'h1 << 45 ) : p ;
      p = a [ 7 ] & b [ 39 ] ? p + ( 60'h1 << 46 ) : p ;
      p = a [ 7 ] & b [ 40 ] ? p + ( 60'h1 << 47 ) : p ;
      p = a [ 7 ] & b [ 41 ] ? p + ( 60'h1 << 48 ) : p ;
      p = a [ 7 ] & b [ 42 ] ? p + ( 60'h1 << 49 ) : p ;
      p = a [ 7 ] & b [ 43 ] ? p + ( 60'h1 << 50 ) : p ;
      p = a [ 7 ] & b [ 44 ] ? p + ( 60'h1 << 51 ) : p ;
      p = a [ 7 ] & b [ 45 ] ? p + ( 60'h1 << 52 ) : p ;
      p = a [ 7 ] & b [ 46 ] ? p + ( 60'h1 << 53 ) : p ;
      p = a [ 7 ] & b [ 47 ] ? p + ( 60'h1 << 54 ) : p ;
      p = a [ 7 ] & b [ 48 ] ? p + ( 60'h1 << 55 ) : p ;
      p = a [ 7 ] & b [ 49 ] ? p + ( 60'h1 << 56 ) : p ;
      p = a [ 7 ] & b [ 50 ] ? p + ( 60'h1 << 57 ) : p ;
      p = a [ 7 ] & b [ 51 ] ? p + ( 60'h1 << 58 ) : p ;
      p = a [ 7 ] & b [ 52 ] ? p + ( 60'h1 << 59 ) : p ;

// Bit by Bit Multiply & Divide + Modulus
// Copyright © 2022 by Gregory Scott Callen
// All Rights Reserved.

      p = a [ 8 ] & b [ 0 ] ? p + ( 60'h1 << 8 ) : p ;
      p = a [ 8 ] & b [ 1 ] ? p + ( 60'h1 << 9 ) : p ;
      p = a [ 8 ] & b [ 2 ] ? p + ( 60'h1 << 10 ) : p ;
      p = a [ 8 ] & b [ 3 ] ? p + ( 60'h1 << 11 ) : p ;
      p = a [ 8 ] & b [ 4 ] ? p + ( 60'h1 << 12 ) : p ;
      p = a [ 8 ] & b [ 5 ] ? p + ( 60'h1 << 13 ) : p ;
      p = a [ 8 ] & b [ 6 ] ? p + ( 60'h1 << 14 ) : p ;
      p = a [ 8 ] & b [ 7 ] ? p + ( 60'h1 << 15 ) : p ;
      p = a [ 8 ] & b [ 8 ] ? p + ( 60'h1 << 16 ) : p ;
      p = a [ 8 ] & b [ 9 ] ? p + ( 60'h1 << 17 ) : p ;
      p = a [ 8 ] & b [ 10 ] ? p + ( 60'h1 << 18 ) : p ;
      p = a [ 8 ] & b [ 11 ] ? p + ( 60'h1 << 19 ) : p ;
      p = a [ 8 ] & b [ 12 ] ? p + ( 60'h1 << 20 ) : p ;
      p = a [ 8 ] & b [ 13 ] ? p + ( 60'h1 << 21 ) : p ;
      p = a [ 8 ] & b [ 14 ] ? p + ( 60'h1 << 22 ) : p ;
      p = a [ 8 ] & b [ 15 ] ? p + ( 60'h1 << 23 ) : p ;
      p = a [ 8 ] & b [ 16 ] ? p + ( 60'h1 << 24 ) : p ;
      p = a [ 8 ] & b [ 17 ] ? p + ( 60'h1 << 25 ) : p ;
      p = a [ 8 ] & b [ 18 ] ? p + ( 60'h1 << 26 ) : p ;
      p = a [ 8 ] & b [ 19 ] ? p + ( 60'h1 << 27 ) : p ;
      p = a [ 8 ] & b [ 20 ] ? p + ( 60'h1 << 28 ) : p ;
      p = a [ 8 ] & b [ 21 ] ? p + ( 60'h1 << 29 ) : p ;
      p = a [ 8 ] & b [ 22 ] ? p + ( 60'h1 << 30 ) : p ;
      p = a [ 8 ] & b [ 23 ] ? p + ( 60'h1 << 31 ) : p ;
      p = a [ 8 ] & b [ 24 ] ? p + ( 60'h1 << 32 ) : p ;
      p = a [ 8 ] & b [ 25 ] ? p + ( 60'h1 << 33 ) : p ;
      p = a [ 8 ] & b [ 26 ] ? p + ( 60'h1 << 34 ) : p ;
      p = a [ 8 ] & b [ 27 ] ? p + ( 60'h1 << 35 ) : p ;
      p = a [ 8 ] & b [ 28 ] ? p + ( 60'h1 << 36 ) : p ;
      p = a [ 8 ] & b [ 29 ] ? p + ( 60'h1 << 37 ) : p ;
      p = a [ 8 ] & b [ 30 ] ? p + ( 60'h1 << 38 ) : p ;
      p = a [ 8 ] & b [ 31 ] ? p + ( 60'h1 << 39 ) : p ;
      p = a [ 8 ] & b [ 32 ] ? p + ( 60'h1 << 40 ) : p ;
      p = a [ 8 ] & b [ 33 ] ? p + ( 60'h1 << 41 ) : p ;
      p = a [ 8 ] & b [ 34 ] ? p + ( 60'h1 << 42 ) : p ;
      p = a [ 8 ] & b [ 35 ] ? p + ( 60'h1 << 43 ) : p ;
      p = a [ 8 ] & b [ 36 ] ? p + ( 60'h1 << 44 ) : p ;
      p = a [ 8 ] & b [ 37 ] ? p + ( 60'h1 << 45 ) : p ;
      p = a [ 8 ] & b [ 38 ] ? p + ( 60'h1 << 46 ) : p ;
      p = a [ 8 ] & b [ 39 ] ? p + ( 60'h1 << 47 ) : p ;
      p = a [ 8 ] & b [ 40 ] ? p + ( 60'h1 << 48 ) : p ;
      p = a [ 8 ] & b [ 41 ] ? p + ( 60'h1 << 49 ) : p ;
      p = a [ 8 ] & b [ 42 ] ? p + ( 60'h1 << 50 ) : p ;
      p = a [ 8 ] & b [ 43 ] ? p + ( 60'h1 << 51 ) : p ;
      p = a [ 8 ] & b [ 44 ] ? p + ( 60'h1 << 52 ) : p ;
      p = a [ 8 ] & b [ 45 ] ? p + ( 60'h1 << 53 ) : p ;
      p = a [ 8 ] & b [ 46 ] ? p + ( 60'h1 << 54 ) : p ;
      p = a [ 8 ] & b [ 47 ] ? p + ( 60'h1 << 55 ) : p ;
      p = a [ 8 ] & b [ 48 ] ? p + ( 60'h1 << 56 ) : p ;
      p = a [ 8 ] & b [ 49 ] ? p + ( 60'h1 << 57 ) : p ;
      p = a [ 8 ] & b [ 50 ] ? p + ( 60'h1 << 58 ) : p ;
      p = a [ 8 ] & b [ 51 ] ? p + ( 60'h1 << 59 ) : p ;

// Bit by Bit Multiply & Divide + Modulus
// Copyright © 2022 by Gregory Scott Callen
// All Rights Reserved.

      p = a [ 9 ] & b [ 0 ] ? p + ( 60'h1 << 9 ) : p ;
      p = a [ 9 ] & b [ 1 ] ? p + ( 60'h1 << 10 ) : p ;
      p = a [ 9 ] & b [ 2 ] ? p + ( 60'h1 << 11 ) : p ;
      p = a [ 9 ] & b [ 3 ] ? p + ( 60'h1 << 12 ) : p ;
      p = a [ 9 ] & b [ 4 ] ? p + ( 60'h1 << 13 ) : p ;
      p = a [ 9 ] & b [ 5 ] ? p + ( 60'h1 << 14 ) : p ;
      p = a [ 9 ] & b [ 6 ] ? p + ( 60'h1 << 15 ) : p ;
      p = a [ 9 ] & b [ 7 ] ? p + ( 60'h1 << 16 ) : p ;
      p = a [ 9 ] & b [ 8 ] ? p + ( 60'h1 << 17 ) : p ;
      p = a [ 9 ] & b [ 9 ] ? p + ( 60'h1 << 18 ) : p ;
      p = a [ 9 ] & b [ 10 ] ? p + ( 60'h1 << 19 ) : p ;
      p = a [ 9 ] & b [ 11 ] ? p + ( 60'h1 << 20 ) : p ;
      p = a [ 9 ] & b [ 12 ] ? p + ( 60'h1 << 21 ) : p ;
      p = a [ 9 ] & b [ 13 ] ? p + ( 60'h1 << 22 ) : p ;
      p = a [ 9 ] & b [ 14 ] ? p + ( 60'h1 << 23 ) : p ;
      p = a [ 9 ] & b [ 15 ] ? p + ( 60'h1 << 24 ) : p ;
      p = a [ 9 ] & b [ 16 ] ? p + ( 60'h1 << 25 ) : p ;
      p = a [ 9 ] & b [ 17 ] ? p + ( 60'h1 << 26 ) : p ;
      p = a [ 9 ] & b [ 18 ] ? p + ( 60'h1 << 27 ) : p ;
      p = a [ 9 ] & b [ 19 ] ? p + ( 60'h1 << 28 ) : p ;
      p = a [ 9 ] & b [ 20 ] ? p + ( 60'h1 << 29 ) : p ;
      p = a [ 9 ] & b [ 21 ] ? p + ( 60'h1 << 30 ) : p ;
      p = a [ 9 ] & b [ 22 ] ? p + ( 60'h1 << 31 ) : p ;
      p = a [ 9 ] & b [ 23 ] ? p + ( 60'h1 << 32 ) : p ;
      p = a [ 9 ] & b [ 24 ] ? p + ( 60'h1 << 33 ) : p ;
      p = a [ 9 ] & b [ 25 ] ? p + ( 60'h1 << 34 ) : p ;
      p = a [ 9 ] & b [ 26 ] ? p + ( 60'h1 << 35 ) : p ;
      p = a [ 9 ] & b [ 27 ] ? p + ( 60'h1 << 36 ) : p ;
      p = a [ 9 ] & b [ 28 ] ? p + ( 60'h1 << 37 ) : p ;
      p = a [ 9 ] & b [ 29 ] ? p + ( 60'h1 << 38 ) : p ;
      p = a [ 9 ] & b [ 30 ] ? p + ( 60'h1 << 39 ) : p ;
      p = a [ 9 ] & b [ 31 ] ? p + ( 60'h1 << 40 ) : p ;
      p = a [ 9 ] & b [ 32 ] ? p + ( 60'h1 << 41 ) : p ;
      p = a [ 9 ] & b [ 33 ] ? p + ( 60'h1 << 42 ) : p ;
      p = a [ 9 ] & b [ 34 ] ? p + ( 60'h1 << 43 ) : p ;
      p = a [ 9 ] & b [ 35 ] ? p + ( 60'h1 << 44 ) : p ;
      p = a [ 9 ] & b [ 36 ] ? p + ( 60'h1 << 45 ) : p ;
      p = a [ 9 ] & b [ 37 ] ? p + ( 60'h1 << 46 ) : p ;
      p = a [ 9 ] & b [ 38 ] ? p + ( 60'h1 << 47 ) : p ;
      p = a [ 9 ] & b [ 39 ] ? p + ( 60'h1 << 48 ) : p ;
      p = a [ 9 ] & b [ 40 ] ? p + ( 60'h1 << 49 ) : p ;
      p = a [ 9 ] & b [ 41 ] ? p + ( 60'h1 << 50 ) : p ;
      p = a [ 9 ] & b [ 42 ] ? p + ( 60'h1 << 51 ) : p ;
      p = a [ 9 ] & b [ 43 ] ? p + ( 60'h1 << 52 ) : p ;
      p = a [ 9 ] & b [ 44 ] ? p + ( 60'h1 << 53 ) : p ;
      p = a [ 9 ] & b [ 45 ] ? p + ( 60'h1 << 54 ) : p ;
      p = a [ 9 ] & b [ 46 ] ? p + ( 60'h1 << 55 ) : p ;
      p = a [ 9 ] & b [ 47 ] ? p + ( 60'h1 << 56 ) : p ;
      p = a [ 9 ] & b [ 48 ] ? p + ( 60'h1 << 57 ) : p ;
      p = a [ 9 ] & b [ 49 ] ? p + ( 60'h1 << 58 ) : p ;
      p = a [ 9 ] & b [ 50 ] ? p + ( 60'h1 << 59 ) : p ;

// Bit by Bit Multiply & Divide + Modulus
// Copyright © 2022 by Gregory Scott Callen
// All Rights Reserved.

      p = a [ 10 ] & b [ 0 ] ? p + ( 60'h1 << 10 ) : p ;
      p = a [ 10 ] & b [ 1 ] ? p + ( 60'h1 << 11 ) : p ;
      p = a [ 10 ] & b [ 2 ] ? p + ( 60'h1 << 12 ) : p ;
      p = a [ 10 ] & b [ 3 ] ? p + ( 60'h1 << 13 ) : p ;
      p = a [ 10 ] & b [ 4 ] ? p + ( 60'h1 << 14 ) : p ;
      p = a [ 10 ] & b [ 5 ] ? p + ( 60'h1 << 15 ) : p ;
      p = a [ 10 ] & b [ 6 ] ? p + ( 60'h1 << 16 ) : p ;
      p = a [ 10 ] & b [ 7 ] ? p + ( 60'h1 << 17 ) : p ;
      p = a [ 10 ] & b [ 8 ] ? p + ( 60'h1 << 18 ) : p ;
      p = a [ 10 ] & b [ 9 ] ? p + ( 60'h1 << 19 ) : p ;
      p = a [ 10 ] & b [ 10 ] ? p + ( 60'h1 << 20 ) : p ;
      p = a [ 10 ] & b [ 11 ] ? p + ( 60'h1 << 21 ) : p ;
      p = a [ 10 ] & b [ 12 ] ? p + ( 60'h1 << 22 ) : p ;
      p = a [ 10 ] & b [ 13 ] ? p + ( 60'h1 << 23 ) : p ;
      p = a [ 10 ] & b [ 14 ] ? p + ( 60'h1 << 24 ) : p ;
      p = a [ 10 ] & b [ 15 ] ? p + ( 60'h1 << 25 ) : p ;
      p = a [ 10 ] & b [ 16 ] ? p + ( 60'h1 << 26 ) : p ;
      p = a [ 10 ] & b [ 17 ] ? p + ( 60'h1 << 27 ) : p ;
      p = a [ 10 ] & b [ 18 ] ? p + ( 60'h1 << 28 ) : p ;
      p = a [ 10 ] & b [ 19 ] ? p + ( 60'h1 << 29 ) : p ;
      p = a [ 10 ] & b [ 20 ] ? p + ( 60'h1 << 30 ) : p ;
      p = a [ 10 ] & b [ 21 ] ? p + ( 60'h1 << 31 ) : p ;
      p = a [ 10 ] & b [ 22 ] ? p + ( 60'h1 << 32 ) : p ;
      p = a [ 10 ] & b [ 23 ] ? p + ( 60'h1 << 33 ) : p ;
      p = a [ 10 ] & b [ 24 ] ? p + ( 60'h1 << 34 ) : p ;
      p = a [ 10 ] & b [ 25 ] ? p + ( 60'h1 << 35 ) : p ;
      p = a [ 10 ] & b [ 26 ] ? p + ( 60'h1 << 36 ) : p ;
      p = a [ 10 ] & b [ 27 ] ? p + ( 60'h1 << 37 ) : p ;
      p = a [ 10 ] & b [ 28 ] ? p + ( 60'h1 << 38 ) : p ;
      p = a [ 10 ] & b [ 29 ] ? p + ( 60'h1 << 39 ) : p ;
      p = a [ 10 ] & b [ 30 ] ? p + ( 60'h1 << 40 ) : p ;
      p = a [ 10 ] & b [ 31 ] ? p + ( 60'h1 << 41 ) : p ;
      p = a [ 10 ] & b [ 32 ] ? p + ( 60'h1 << 42 ) : p ;
      p = a [ 10 ] & b [ 33 ] ? p + ( 60'h1 << 43 ) : p ;
      p = a [ 10 ] & b [ 34 ] ? p + ( 60'h1 << 44 ) : p ;
      p = a [ 10 ] & b [ 35 ] ? p + ( 60'h1 << 45 ) : p ;
      p = a [ 10 ] & b [ 36 ] ? p + ( 60'h1 << 46 ) : p ;
      p = a [ 10 ] & b [ 37 ] ? p + ( 60'h1 << 47 ) : p ;
      p = a [ 10 ] & b [ 38 ] ? p + ( 60'h1 << 48 ) : p ;
      p = a [ 10 ] & b [ 39 ] ? p + ( 60'h1 << 49 ) : p ;
      p = a [ 10 ] & b [ 40 ] ? p + ( 60'h1 << 50 ) : p ;
      p = a [ 10 ] & b [ 41 ] ? p + ( 60'h1 << 51 ) : p ;
      p = a [ 10 ] & b [ 42 ] ? p + ( 60'h1 << 52 ) : p ;
      p = a [ 10 ] & b [ 43 ] ? p + ( 60'h1 << 53 ) : p ;
      p = a [ 10 ] & b [ 44 ] ? p + ( 60'h1 << 54 ) : p ;
      p = a [ 10 ] & b [ 45 ] ? p + ( 60'h1 << 55 ) : p ;
      p = a [ 10 ] & b [ 46 ] ? p + ( 60'h1 << 56 ) : p ;
      p = a [ 10 ] & b [ 47 ] ? p + ( 60'h1 << 57 ) : p ;
      p = a [ 10 ] & b [ 48 ] ? p + ( 60'h1 << 58 ) : p ;
      p = a [ 10 ] & b [ 49 ] ? p + ( 60'h1 << 59 ) : p ;

// Bit by Bit Multiply & Divide + Modulus
// Copyright © 2022 by Gregory Scott Callen
// All Rights Reserved.

      p = a [ 11 ] & b [ 0 ] ? p + ( 60'h1 << 11 ) : p ;
      p = a [ 11 ] & b [ 1 ] ? p + ( 60'h1 << 12 ) : p ;
      p = a [ 11 ] & b [ 2 ] ? p + ( 60'h1 << 13 ) : p ;
      p = a [ 11 ] & b [ 3 ] ? p + ( 60'h1 << 14 ) : p ;
      p = a [ 11 ] & b [ 4 ] ? p + ( 60'h1 << 15 ) : p ;
      p = a [ 11 ] & b [ 5 ] ? p + ( 60'h1 << 16 ) : p ;
      p = a [ 11 ] & b [ 6 ] ? p + ( 60'h1 << 17 ) : p ;
      p = a [ 11 ] & b [ 7 ] ? p + ( 60'h1 << 18 ) : p ;
      p = a [ 11 ] & b [ 8 ] ? p + ( 60'h1 << 19 ) : p ;
      p = a [ 11 ] & b [ 9 ] ? p + ( 60'h1 << 20 ) : p ;
      p = a [ 11 ] & b [ 10 ] ? p + ( 60'h1 << 21 ) : p ;
      p = a [ 11 ] & b [ 11 ] ? p + ( 60'h1 << 22 ) : p ;
      p = a [ 11 ] & b [ 12 ] ? p + ( 60'h1 << 23 ) : p ;
      p = a [ 11 ] & b [ 13 ] ? p + ( 60'h1 << 24 ) : p ;
      p = a [ 11 ] & b [ 14 ] ? p + ( 60'h1 << 25 ) : p ;
      p = a [ 11 ] & b [ 15 ] ? p + ( 60'h1 << 26 ) : p ;
      p = a [ 11 ] & b [ 16 ] ? p + ( 60'h1 << 27 ) : p ;
      p = a [ 11 ] & b [ 17 ] ? p + ( 60'h1 << 28 ) : p ;
      p = a [ 11 ] & b [ 18 ] ? p + ( 60'h1 << 29 ) : p ;
      p = a [ 11 ] & b [ 19 ] ? p + ( 60'h1 << 30 ) : p ;
      p = a [ 11 ] & b [ 20 ] ? p + ( 60'h1 << 31 ) : p ;
      p = a [ 11 ] & b [ 21 ] ? p + ( 60'h1 << 32 ) : p ;
      p = a [ 11 ] & b [ 22 ] ? p + ( 60'h1 << 33 ) : p ;
      p = a [ 11 ] & b [ 23 ] ? p + ( 60'h1 << 34 ) : p ;
      p = a [ 11 ] & b [ 24 ] ? p + ( 60'h1 << 35 ) : p ;
      p = a [ 11 ] & b [ 25 ] ? p + ( 60'h1 << 36 ) : p ;
      p = a [ 11 ] & b [ 26 ] ? p + ( 60'h1 << 37 ) : p ;
      p = a [ 11 ] & b [ 27 ] ? p + ( 60'h1 << 38 ) : p ;
      p = a [ 11 ] & b [ 28 ] ? p + ( 60'h1 << 39 ) : p ;
      p = a [ 11 ] & b [ 29 ] ? p + ( 60'h1 << 40 ) : p ;
      p = a [ 11 ] & b [ 30 ] ? p + ( 60'h1 << 41 ) : p ;
      p = a [ 11 ] & b [ 31 ] ? p + ( 60'h1 << 42 ) : p ;
      p = a [ 11 ] & b [ 32 ] ? p + ( 60'h1 << 43 ) : p ;
      p = a [ 11 ] & b [ 33 ] ? p + ( 60'h1 << 44 ) : p ;
      p = a [ 11 ] & b [ 34 ] ? p + ( 60'h1 << 45 ) : p ;
      p = a [ 11 ] & b [ 35 ] ? p + ( 60'h1 << 46 ) : p ;
      p = a [ 11 ] & b [ 36 ] ? p + ( 60'h1 << 47 ) : p ;
      p = a [ 11 ] & b [ 37 ] ? p + ( 60'h1 << 48 ) : p ;
      p = a [ 11 ] & b [ 38 ] ? p + ( 60'h1 << 49 ) : p ;
      p = a [ 11 ] & b [ 39 ] ? p + ( 60'h1 << 50 ) : p ;
      p = a [ 11 ] & b [ 40 ] ? p + ( 60'h1 << 51 ) : p ;
      p = a [ 11 ] & b [ 41 ] ? p + ( 60'h1 << 52 ) : p ;
      p = a [ 11 ] & b [ 42 ] ? p + ( 60'h1 << 53 ) : p ;
      p = a [ 11 ] & b [ 43 ] ? p + ( 60'h1 << 54 ) : p ;
      p = a [ 11 ] & b [ 44 ] ? p + ( 60'h1 << 55 ) : p ;
      p = a [ 11 ] & b [ 45 ] ? p + ( 60'h1 << 56 ) : p ;
      p = a [ 11 ] & b [ 46 ] ? p + ( 60'h1 << 57 ) : p ;
      p = a [ 11 ] & b [ 47 ] ? p + ( 60'h1 << 58 ) : p ;
      p = a [ 11 ] & b [ 48 ] ? p + ( 60'h1 << 59 ) : p ;

// Bit by Bit Multiply & Divide + Modulus
// Copyright © 2022 by Gregory Scott Callen
// All Rights Reserved.

      p = a [ 12 ] & b [ 0 ] ? p + ( 60'h1 << 12 ) : p ;
      p = a [ 12 ] & b [ 1 ] ? p + ( 60'h1 << 13 ) : p ;
      p = a [ 12 ] & b [ 2 ] ? p + ( 60'h1 << 14 ) : p ;
      p = a [ 12 ] & b [ 3 ] ? p + ( 60'h1 << 15 ) : p ;
      p = a [ 12 ] & b [ 4 ] ? p + ( 60'h1 << 16 ) : p ;
      p = a [ 12 ] & b [ 5 ] ? p + ( 60'h1 << 17 ) : p ;
      p = a [ 12 ] & b [ 6 ] ? p + ( 60'h1 << 18 ) : p ;
      p = a [ 12 ] & b [ 7 ] ? p + ( 60'h1 << 19 ) : p ;
      p = a [ 12 ] & b [ 8 ] ? p + ( 60'h1 << 20 ) : p ;
      p = a [ 12 ] & b [ 9 ] ? p + ( 60'h1 << 21 ) : p ;
      p = a [ 12 ] & b [ 10 ] ? p + ( 60'h1 << 22 ) : p ;
      p = a [ 12 ] & b [ 11 ] ? p + ( 60'h1 << 23 ) : p ;
      p = a [ 12 ] & b [ 12 ] ? p + ( 60'h1 << 24 ) : p ;
      p = a [ 12 ] & b [ 13 ] ? p + ( 60'h1 << 25 ) : p ;
      p = a [ 12 ] & b [ 14 ] ? p + ( 60'h1 << 26 ) : p ;
      p = a [ 12 ] & b [ 15 ] ? p + ( 60'h1 << 27 ) : p ;
      p = a [ 12 ] & b [ 16 ] ? p + ( 60'h1 << 28 ) : p ;
      p = a [ 12 ] & b [ 17 ] ? p + ( 60'h1 << 29 ) : p ;
      p = a [ 12 ] & b [ 18 ] ? p + ( 60'h1 << 30 ) : p ;
      p = a [ 12 ] & b [ 19 ] ? p + ( 60'h1 << 31 ) : p ;
      p = a [ 12 ] & b [ 20 ] ? p + ( 60'h1 << 32 ) : p ;
      p = a [ 12 ] & b [ 21 ] ? p + ( 60'h1 << 33 ) : p ;
      p = a [ 12 ] & b [ 22 ] ? p + ( 60'h1 << 34 ) : p ;
      p = a [ 12 ] & b [ 23 ] ? p + ( 60'h1 << 35 ) : p ;
      p = a [ 12 ] & b [ 24 ] ? p + ( 60'h1 << 36 ) : p ;
      p = a [ 12 ] & b [ 25 ] ? p + ( 60'h1 << 37 ) : p ;
      p = a [ 12 ] & b [ 26 ] ? p + ( 60'h1 << 38 ) : p ;
      p = a [ 12 ] & b [ 27 ] ? p + ( 60'h1 << 39 ) : p ;
      p = a [ 12 ] & b [ 28 ] ? p + ( 60'h1 << 40 ) : p ;
      p = a [ 12 ] & b [ 29 ] ? p + ( 60'h1 << 41 ) : p ;
      p = a [ 12 ] & b [ 30 ] ? p + ( 60'h1 << 42 ) : p ;
      p = a [ 12 ] & b [ 31 ] ? p + ( 60'h1 << 43 ) : p ;
      p = a [ 12 ] & b [ 32 ] ? p + ( 60'h1 << 44 ) : p ;
      p = a [ 12 ] & b [ 33 ] ? p + ( 60'h1 << 45 ) : p ;
      p = a [ 12 ] & b [ 34 ] ? p + ( 60'h1 << 46 ) : p ;
      p = a [ 12 ] & b [ 35 ] ? p + ( 60'h1 << 47 ) : p ;
      p = a [ 12 ] & b [ 36 ] ? p + ( 60'h1 << 48 ) : p ;
      p = a [ 12 ] & b [ 37 ] ? p + ( 60'h1 << 49 ) : p ;
      p = a [ 12 ] & b [ 38 ] ? p + ( 60'h1 << 50 ) : p ;
      p = a [ 12 ] & b [ 39 ] ? p + ( 60'h1 << 51 ) : p ;
      p = a [ 12 ] & b [ 40 ] ? p + ( 60'h1 << 52 ) : p ;
      p = a [ 12 ] & b [ 41 ] ? p + ( 60'h1 << 53 ) : p ;
      p = a [ 12 ] & b [ 42 ] ? p + ( 60'h1 << 54 ) : p ;
      p = a [ 12 ] & b [ 43 ] ? p + ( 60'h1 << 55 ) : p ;
      p = a [ 12 ] & b [ 44 ] ? p + ( 60'h1 << 56 ) : p ;
      p = a [ 12 ] & b [ 45 ] ? p + ( 60'h1 << 57 ) : p ;
      p = a [ 12 ] & b [ 46 ] ? p + ( 60'h1 << 58 ) : p ;
      p = a [ 12 ] & b [ 47 ] ? p + ( 60'h1 << 59 ) : p ;

// Bit by Bit Multiply & Divide + Modulus
// Copyright © 2022 by Gregory Scott Callen
// All Rights Reserved.

      p = a [ 13 ] & b [ 0 ] ? p + ( 60'h1 << 13 ) : p ;
      p = a [ 13 ] & b [ 1 ] ? p + ( 60'h1 << 14 ) : p ;
      p = a [ 13 ] & b [ 2 ] ? p + ( 60'h1 << 15 ) : p ;
      p = a [ 13 ] & b [ 3 ] ? p + ( 60'h1 << 16 ) : p ;
      p = a [ 13 ] & b [ 4 ] ? p + ( 60'h1 << 17 ) : p ;
      p = a [ 13 ] & b [ 5 ] ? p + ( 60'h1 << 18 ) : p ;
      p = a [ 13 ] & b [ 6 ] ? p + ( 60'h1 << 19 ) : p ;
      p = a [ 13 ] & b [ 7 ] ? p + ( 60'h1 << 20 ) : p ;
      p = a [ 13 ] & b [ 8 ] ? p + ( 60'h1 << 21 ) : p ;
      p = a [ 13 ] & b [ 9 ] ? p + ( 60'h1 << 22 ) : p ;
      p = a [ 13 ] & b [ 10 ] ? p + ( 60'h1 << 23 ) : p ;
      p = a [ 13 ] & b [ 11 ] ? p + ( 60'h1 << 24 ) : p ;
      p = a [ 13 ] & b [ 12 ] ? p + ( 60'h1 << 25 ) : p ;
      p = a [ 13 ] & b [ 13 ] ? p + ( 60'h1 << 26 ) : p ;
      p = a [ 13 ] & b [ 14 ] ? p + ( 60'h1 << 27 ) : p ;
      p = a [ 13 ] & b [ 15 ] ? p + ( 60'h1 << 28 ) : p ;
      p = a [ 13 ] & b [ 16 ] ? p + ( 60'h1 << 29 ) : p ;
      p = a [ 13 ] & b [ 17 ] ? p + ( 60'h1 << 30 ) : p ;
      p = a [ 13 ] & b [ 18 ] ? p + ( 60'h1 << 31 ) : p ;
      p = a [ 13 ] & b [ 19 ] ? p + ( 60'h1 << 32 ) : p ;
      p = a [ 13 ] & b [ 20 ] ? p + ( 60'h1 << 33 ) : p ;
      p = a [ 13 ] & b [ 21 ] ? p + ( 60'h1 << 34 ) : p ;
      p = a [ 13 ] & b [ 22 ] ? p + ( 60'h1 << 35 ) : p ;
      p = a [ 13 ] & b [ 23 ] ? p + ( 60'h1 << 36 ) : p ;
      p = a [ 13 ] & b [ 24 ] ? p + ( 60'h1 << 37 ) : p ;
      p = a [ 13 ] & b [ 25 ] ? p + ( 60'h1 << 38 ) : p ;
      p = a [ 13 ] & b [ 26 ] ? p + ( 60'h1 << 39 ) : p ;
      p = a [ 13 ] & b [ 27 ] ? p + ( 60'h1 << 40 ) : p ;
      p = a [ 13 ] & b [ 28 ] ? p + ( 60'h1 << 41 ) : p ;
      p = a [ 13 ] & b [ 29 ] ? p + ( 60'h1 << 42 ) : p ;
      p = a [ 13 ] & b [ 30 ] ? p + ( 60'h1 << 43 ) : p ;
      p = a [ 13 ] & b [ 31 ] ? p + ( 60'h1 << 44 ) : p ;
      p = a [ 13 ] & b [ 32 ] ? p + ( 60'h1 << 45 ) : p ;
      p = a [ 13 ] & b [ 33 ] ? p + ( 60'h1 << 46 ) : p ;
      p = a [ 13 ] & b [ 34 ] ? p + ( 60'h1 << 47 ) : p ;
      p = a [ 13 ] & b [ 35 ] ? p + ( 60'h1 << 48 ) : p ;
      p = a [ 13 ] & b [ 36 ] ? p + ( 60'h1 << 49 ) : p ;
      p = a [ 13 ] & b [ 37 ] ? p + ( 60'h1 << 50 ) : p ;
      p = a [ 13 ] & b [ 38 ] ? p + ( 60'h1 << 51 ) : p ;
      p = a [ 13 ] & b [ 39 ] ? p + ( 60'h1 << 52 ) : p ;
      p = a [ 13 ] & b [ 40 ] ? p + ( 60'h1 << 53 ) : p ;
      p = a [ 13 ] & b [ 41 ] ? p + ( 60'h1 << 54 ) : p ;
      p = a [ 13 ] & b [ 42 ] ? p + ( 60'h1 << 55 ) : p ;
      p = a [ 13 ] & b [ 43 ] ? p + ( 60'h1 << 56 ) : p ;
      p = a [ 13 ] & b [ 44 ] ? p + ( 60'h1 << 57 ) : p ;
      p = a [ 13 ] & b [ 45 ] ? p + ( 60'h1 << 58 ) : p ;
      p = a [ 13 ] & b [ 46 ] ? p + ( 60'h1 << 59 ) : p ;

// Bit by Bit Multiply & Divide + Modulus
// Copyright © 2022 by Gregory Scott Callen
// All Rights Reserved.

      p = a [ 14 ] & b [ 0 ] ? p + ( 60'h1 << 14 ) : p ;
      p = a [ 14 ] & b [ 1 ] ? p + ( 60'h1 << 15 ) : p ;
      p = a [ 14 ] & b [ 2 ] ? p + ( 60'h1 << 16 ) : p ;
      p = a [ 14 ] & b [ 3 ] ? p + ( 60'h1 << 17 ) : p ;
      p = a [ 14 ] & b [ 4 ] ? p + ( 60'h1 << 18 ) : p ;
      p = a [ 14 ] & b [ 5 ] ? p + ( 60'h1 << 19 ) : p ;
      p = a [ 14 ] & b [ 6 ] ? p + ( 60'h1 << 20 ) : p ;
      p = a [ 14 ] & b [ 7 ] ? p + ( 60'h1 << 21 ) : p ;
      p = a [ 14 ] & b [ 8 ] ? p + ( 60'h1 << 22 ) : p ;
      p = a [ 14 ] & b [ 9 ] ? p + ( 60'h1 << 23 ) : p ;
      p = a [ 14 ] & b [ 10 ] ? p + ( 60'h1 << 24 ) : p ;
      p = a [ 14 ] & b [ 11 ] ? p + ( 60'h1 << 25 ) : p ;
      p = a [ 14 ] & b [ 12 ] ? p + ( 60'h1 << 26 ) : p ;
      p = a [ 14 ] & b [ 13 ] ? p + ( 60'h1 << 27 ) : p ;
      p = a [ 14 ] & b [ 14 ] ? p + ( 60'h1 << 28 ) : p ;
      p = a [ 14 ] & b [ 15 ] ? p + ( 60'h1 << 29 ) : p ;
      p = a [ 14 ] & b [ 16 ] ? p + ( 60'h1 << 30 ) : p ;
      p = a [ 14 ] & b [ 17 ] ? p + ( 60'h1 << 31 ) : p ;
      p = a [ 14 ] & b [ 18 ] ? p + ( 60'h1 << 32 ) : p ;
      p = a [ 14 ] & b [ 19 ] ? p + ( 60'h1 << 33 ) : p ;
      p = a [ 14 ] & b [ 20 ] ? p + ( 60'h1 << 34 ) : p ;
      p = a [ 14 ] & b [ 21 ] ? p + ( 60'h1 << 35 ) : p ;
      p = a [ 14 ] & b [ 22 ] ? p + ( 60'h1 << 36 ) : p ;
      p = a [ 14 ] & b [ 23 ] ? p + ( 60'h1 << 37 ) : p ;
      p = a [ 14 ] & b [ 24 ] ? p + ( 60'h1 << 38 ) : p ;
      p = a [ 14 ] & b [ 25 ] ? p + ( 60'h1 << 39 ) : p ;
      p = a [ 14 ] & b [ 26 ] ? p + ( 60'h1 << 40 ) : p ;
      p = a [ 14 ] & b [ 27 ] ? p + ( 60'h1 << 41 ) : p ;
      p = a [ 14 ] & b [ 28 ] ? p + ( 60'h1 << 42 ) : p ;
      p = a [ 14 ] & b [ 29 ] ? p + ( 60'h1 << 43 ) : p ;
      p = a [ 14 ] & b [ 30 ] ? p + ( 60'h1 << 44 ) : p ;
      p = a [ 14 ] & b [ 31 ] ? p + ( 60'h1 << 45 ) : p ;
      p = a [ 14 ] & b [ 32 ] ? p + ( 60'h1 << 46 ) : p ;
      p = a [ 14 ] & b [ 33 ] ? p + ( 60'h1 << 47 ) : p ;
      p = a [ 14 ] & b [ 34 ] ? p + ( 60'h1 << 48 ) : p ;
      p = a [ 14 ] & b [ 35 ] ? p + ( 60'h1 << 49 ) : p ;
      p = a [ 14 ] & b [ 36 ] ? p + ( 60'h1 << 50 ) : p ;
      p = a [ 14 ] & b [ 37 ] ? p + ( 60'h1 << 51 ) : p ;
      p = a [ 14 ] & b [ 38 ] ? p + ( 60'h1 << 52 ) : p ;
      p = a [ 14 ] & b [ 39 ] ? p + ( 60'h1 << 53 ) : p ;
      p = a [ 14 ] & b [ 40 ] ? p + ( 60'h1 << 54 ) : p ;
      p = a [ 14 ] & b [ 41 ] ? p + ( 60'h1 << 55 ) : p ;
      p = a [ 14 ] & b [ 42 ] ? p + ( 60'h1 << 56 ) : p ;
      p = a [ 14 ] & b [ 43 ] ? p + ( 60'h1 << 57 ) : p ;
      p = a [ 14 ] & b [ 44 ] ? p + ( 60'h1 << 58 ) : p ;
      p = a [ 14 ] & b [ 45 ] ? p + ( 60'h1 << 59 ) : p ;

// Bit by Bit Multiply & Divide + Modulus
// Copyright © 2022 by Gregory Scott Callen
// All Rights Reserved.

      p = a [ 15 ] & b [ 0 ] ? p + ( 60'h1 << 15 ) : p ;
      p = a [ 15 ] & b [ 1 ] ? p + ( 60'h1 << 16 ) : p ;
      p = a [ 15 ] & b [ 2 ] ? p + ( 60'h1 << 17 ) : p ;
      p = a [ 15 ] & b [ 3 ] ? p + ( 60'h1 << 18 ) : p ;
      p = a [ 15 ] & b [ 4 ] ? p + ( 60'h1 << 19 ) : p ;
      p = a [ 15 ] & b [ 5 ] ? p + ( 60'h1 << 20 ) : p ;
      p = a [ 15 ] & b [ 6 ] ? p + ( 60'h1 << 21 ) : p ;
      p = a [ 15 ] & b [ 7 ] ? p + ( 60'h1 << 22 ) : p ;
      p = a [ 15 ] & b [ 8 ] ? p + ( 60'h1 << 23 ) : p ;
      p = a [ 15 ] & b [ 9 ] ? p + ( 60'h1 << 24 ) : p ;
      p = a [ 15 ] & b [ 10 ] ? p + ( 60'h1 << 25 ) : p ;
      p = a [ 15 ] & b [ 11 ] ? p + ( 60'h1 << 26 ) : p ;
      p = a [ 15 ] & b [ 12 ] ? p + ( 60'h1 << 27 ) : p ;
      p = a [ 15 ] & b [ 13 ] ? p + ( 60'h1 << 28 ) : p ;
      p = a [ 15 ] & b [ 14 ] ? p + ( 60'h1 << 29 ) : p ;
      p = a [ 15 ] & b [ 15 ] ? p + ( 60'h1 << 30 ) : p ;
      p = a [ 15 ] & b [ 16 ] ? p + ( 60'h1 << 31 ) : p ;
      p = a [ 15 ] & b [ 17 ] ? p + ( 60'h1 << 32 ) : p ;
      p = a [ 15 ] & b [ 18 ] ? p + ( 60'h1 << 33 ) : p ;
      p = a [ 15 ] & b [ 19 ] ? p + ( 60'h1 << 34 ) : p ;
      p = a [ 15 ] & b [ 20 ] ? p + ( 60'h1 << 35 ) : p ;
      p = a [ 15 ] & b [ 21 ] ? p + ( 60'h1 << 36 ) : p ;
      p = a [ 15 ] & b [ 22 ] ? p + ( 60'h1 << 37 ) : p ;
      p = a [ 15 ] & b [ 23 ] ? p + ( 60'h1 << 38 ) : p ;
      p = a [ 15 ] & b [ 24 ] ? p + ( 60'h1 << 39 ) : p ;
      p = a [ 15 ] & b [ 25 ] ? p + ( 60'h1 << 40 ) : p ;
      p = a [ 15 ] & b [ 26 ] ? p + ( 60'h1 << 41 ) : p ;
      p = a [ 15 ] & b [ 27 ] ? p + ( 60'h1 << 42 ) : p ;
      p = a [ 15 ] & b [ 28 ] ? p + ( 60'h1 << 43 ) : p ;
      p = a [ 15 ] & b [ 29 ] ? p + ( 60'h1 << 44 ) : p ;
      p = a [ 15 ] & b [ 30 ] ? p + ( 60'h1 << 45 ) : p ;
      p = a [ 15 ] & b [ 31 ] ? p + ( 60'h1 << 46 ) : p ;
      p = a [ 15 ] & b [ 32 ] ? p + ( 60'h1 << 47 ) : p ;
      p = a [ 15 ] & b [ 33 ] ? p + ( 60'h1 << 48 ) : p ;
      p = a [ 15 ] & b [ 34 ] ? p + ( 60'h1 << 49 ) : p ;
      p = a [ 15 ] & b [ 35 ] ? p + ( 60'h1 << 50 ) : p ;
      p = a [ 15 ] & b [ 36 ] ? p + ( 60'h1 << 51 ) : p ;
      p = a [ 15 ] & b [ 37 ] ? p + ( 60'h1 << 52 ) : p ;
      p = a [ 15 ] & b [ 38 ] ? p + ( 60'h1 << 53 ) : p ;
      p = a [ 15 ] & b [ 39 ] ? p + ( 60'h1 << 54 ) : p ;
      p = a [ 15 ] & b [ 40 ] ? p + ( 60'h1 << 55 ) : p ;
      p = a [ 15 ] & b [ 41 ] ? p + ( 60'h1 << 56 ) : p ;
      p = a [ 15 ] & b [ 42 ] ? p + ( 60'h1 << 57 ) : p ;
      p = a [ 15 ] & b [ 43 ] ? p + ( 60'h1 << 58 ) : p ;
      p = a [ 15 ] & b [ 44 ] ? p + ( 60'h1 << 59 ) : p ;

// Bit by Bit Multiply & Divide + Modulus
// Copyright © 2022 by Gregory Scott Callen
// All Rights Reserved.

      p = a [ 16 ] & b [ 0 ] ? p + ( 60'h1 << 16 ) : p ;
      p = a [ 16 ] & b [ 1 ] ? p + ( 60'h1 << 17 ) : p ;
      p = a [ 16 ] & b [ 2 ] ? p + ( 60'h1 << 18 ) : p ;
      p = a [ 16 ] & b [ 3 ] ? p + ( 60'h1 << 19 ) : p ;
      p = a [ 16 ] & b [ 4 ] ? p + ( 60'h1 << 20 ) : p ;
      p = a [ 16 ] & b [ 5 ] ? p + ( 60'h1 << 21 ) : p ;
      p = a [ 16 ] & b [ 6 ] ? p + ( 60'h1 << 22 ) : p ;
      p = a [ 16 ] & b [ 7 ] ? p + ( 60'h1 << 23 ) : p ;
      p = a [ 16 ] & b [ 8 ] ? p + ( 60'h1 << 24 ) : p ;
      p = a [ 16 ] & b [ 9 ] ? p + ( 60'h1 << 25 ) : p ;
      p = a [ 16 ] & b [ 10 ] ? p + ( 60'h1 << 26 ) : p ;
      p = a [ 16 ] & b [ 11 ] ? p + ( 60'h1 << 27 ) : p ;
      p = a [ 16 ] & b [ 12 ] ? p + ( 60'h1 << 28 ) : p ;
      p = a [ 16 ] & b [ 13 ] ? p + ( 60'h1 << 29 ) : p ;
      p = a [ 16 ] & b [ 14 ] ? p + ( 60'h1 << 30 ) : p ;
      p = a [ 16 ] & b [ 15 ] ? p + ( 60'h1 << 31 ) : p ;
      p = a [ 16 ] & b [ 16 ] ? p + ( 60'h1 << 32 ) : p ;
      p = a [ 16 ] & b [ 17 ] ? p + ( 60'h1 << 33 ) : p ;
      p = a [ 16 ] & b [ 18 ] ? p + ( 60'h1 << 34 ) : p ;
      p = a [ 16 ] & b [ 19 ] ? p + ( 60'h1 << 35 ) : p ;
      p = a [ 16 ] & b [ 20 ] ? p + ( 60'h1 << 36 ) : p ;
      p = a [ 16 ] & b [ 21 ] ? p + ( 60'h1 << 37 ) : p ;
      p = a [ 16 ] & b [ 22 ] ? p + ( 60'h1 << 38 ) : p ;
      p = a [ 16 ] & b [ 23 ] ? p + ( 60'h1 << 39 ) : p ;
      p = a [ 16 ] & b [ 24 ] ? p + ( 60'h1 << 40 ) : p ;
      p = a [ 16 ] & b [ 25 ] ? p + ( 60'h1 << 41 ) : p ;
      p = a [ 16 ] & b [ 26 ] ? p + ( 60'h1 << 42 ) : p ;
      p = a [ 16 ] & b [ 27 ] ? p + ( 60'h1 << 43 ) : p ;
      p = a [ 16 ] & b [ 28 ] ? p + ( 60'h1 << 44 ) : p ;
      p = a [ 16 ] & b [ 29 ] ? p + ( 60'h1 << 45 ) : p ;
      p = a [ 16 ] & b [ 30 ] ? p + ( 60'h1 << 46 ) : p ;
      p = a [ 16 ] & b [ 31 ] ? p + ( 60'h1 << 47 ) : p ;
      p = a [ 16 ] & b [ 32 ] ? p + ( 60'h1 << 48 ) : p ;
      p = a [ 16 ] & b [ 33 ] ? p + ( 60'h1 << 49 ) : p ;
      p = a [ 16 ] & b [ 34 ] ? p + ( 60'h1 << 50 ) : p ;
      p = a [ 16 ] & b [ 35 ] ? p + ( 60'h1 << 51 ) : p ;
      p = a [ 16 ] & b [ 36 ] ? p + ( 60'h1 << 52 ) : p ;
      p = a [ 16 ] & b [ 37 ] ? p + ( 60'h1 << 53 ) : p ;
      p = a [ 16 ] & b [ 38 ] ? p + ( 60'h1 << 54 ) : p ;
      p = a [ 16 ] & b [ 39 ] ? p + ( 60'h1 << 55 ) : p ;
      p = a [ 16 ] & b [ 40 ] ? p + ( 60'h1 << 56 ) : p ;
      p = a [ 16 ] & b [ 41 ] ? p + ( 60'h1 << 57 ) : p ;
      p = a [ 16 ] & b [ 42 ] ? p + ( 60'h1 << 58 ) : p ;
      p = a [ 16 ] & b [ 43 ] ? p + ( 60'h1 << 59 ) : p ;

// Bit by Bit Multiply & Divide + Modulus
// Copyright © 2022 by Gregory Scott Callen
// All Rights Reserved.

      p = a [ 17 ] & b [ 0 ] ? p + ( 60'h1 << 17 ) : p ;
      p = a [ 17 ] & b [ 1 ] ? p + ( 60'h1 << 18 ) : p ;
      p = a [ 17 ] & b [ 2 ] ? p + ( 60'h1 << 19 ) : p ;
      p = a [ 17 ] & b [ 3 ] ? p + ( 60'h1 << 20 ) : p ;
      p = a [ 17 ] & b [ 4 ] ? p + ( 60'h1 << 21 ) : p ;
      p = a [ 17 ] & b [ 5 ] ? p + ( 60'h1 << 22 ) : p ;
      p = a [ 17 ] & b [ 6 ] ? p + ( 60'h1 << 23 ) : p ;
      p = a [ 17 ] & b [ 7 ] ? p + ( 60'h1 << 24 ) : p ;
      p = a [ 17 ] & b [ 8 ] ? p + ( 60'h1 << 25 ) : p ;
      p = a [ 17 ] & b [ 9 ] ? p + ( 60'h1 << 26 ) : p ;
      p = a [ 17 ] & b [ 10 ] ? p + ( 60'h1 << 27 ) : p ;
      p = a [ 17 ] & b [ 11 ] ? p + ( 60'h1 << 28 ) : p ;
      p = a [ 17 ] & b [ 12 ] ? p + ( 60'h1 << 29 ) : p ;
      p = a [ 17 ] & b [ 13 ] ? p + ( 60'h1 << 30 ) : p ;
      p = a [ 17 ] & b [ 14 ] ? p + ( 60'h1 << 31 ) : p ;
      p = a [ 17 ] & b [ 15 ] ? p + ( 60'h1 << 32 ) : p ;
      p = a [ 17 ] & b [ 16 ] ? p + ( 60'h1 << 33 ) : p ;
      p = a [ 17 ] & b [ 17 ] ? p + ( 60'h1 << 34 ) : p ;
      p = a [ 17 ] & b [ 18 ] ? p + ( 60'h1 << 35 ) : p ;
      p = a [ 17 ] & b [ 19 ] ? p + ( 60'h1 << 36 ) : p ;
      p = a [ 17 ] & b [ 20 ] ? p + ( 60'h1 << 37 ) : p ;
      p = a [ 17 ] & b [ 21 ] ? p + ( 60'h1 << 38 ) : p ;
      p = a [ 17 ] & b [ 22 ] ? p + ( 60'h1 << 39 ) : p ;
      p = a [ 17 ] & b [ 23 ] ? p + ( 60'h1 << 40 ) : p ;
      p = a [ 17 ] & b [ 24 ] ? p + ( 60'h1 << 41 ) : p ;
      p = a [ 17 ] & b [ 25 ] ? p + ( 60'h1 << 42 ) : p ;
      p = a [ 17 ] & b [ 26 ] ? p + ( 60'h1 << 43 ) : p ;
      p = a [ 17 ] & b [ 27 ] ? p + ( 60'h1 << 44 ) : p ;
      p = a [ 17 ] & b [ 28 ] ? p + ( 60'h1 << 45 ) : p ;
      p = a [ 17 ] & b [ 29 ] ? p + ( 60'h1 << 46 ) : p ;
      p = a [ 17 ] & b [ 30 ] ? p + ( 60'h1 << 47 ) : p ;
      p = a [ 17 ] & b [ 31 ] ? p + ( 60'h1 << 48 ) : p ;
      p = a [ 17 ] & b [ 32 ] ? p + ( 60'h1 << 49 ) : p ;
      p = a [ 17 ] & b [ 33 ] ? p + ( 60'h1 << 50 ) : p ;
      p = a [ 17 ] & b [ 34 ] ? p + ( 60'h1 << 51 ) : p ;
      p = a [ 17 ] & b [ 35 ] ? p + ( 60'h1 << 52 ) : p ;
      p = a [ 17 ] & b [ 36 ] ? p + ( 60'h1 << 53 ) : p ;
      p = a [ 17 ] & b [ 37 ] ? p + ( 60'h1 << 54 ) : p ;
      p = a [ 17 ] & b [ 38 ] ? p + ( 60'h1 << 55 ) : p ;
      p = a [ 17 ] & b [ 39 ] ? p + ( 60'h1 << 56 ) : p ;
      p = a [ 17 ] & b [ 40 ] ? p + ( 60'h1 << 57 ) : p ;
      p = a [ 17 ] & b [ 41 ] ? p + ( 60'h1 << 58 ) : p ;
      p = a [ 17 ] & b [ 42 ] ? p + ( 60'h1 << 59 ) : p ;

// Bit by Bit Multiply & Divide + Modulus
// Copyright © 2022 by Gregory Scott Callen
// All Rights Reserved.

      p = a [ 18 ] & b [ 0 ] ? p + ( 60'h1 << 18 ) : p ;
      p = a [ 18 ] & b [ 1 ] ? p + ( 60'h1 << 19 ) : p ;
      p = a [ 18 ] & b [ 2 ] ? p + ( 60'h1 << 20 ) : p ;
      p = a [ 18 ] & b [ 3 ] ? p + ( 60'h1 << 21 ) : p ;
      p = a [ 18 ] & b [ 4 ] ? p + ( 60'h1 << 22 ) : p ;
      p = a [ 18 ] & b [ 5 ] ? p + ( 60'h1 << 23 ) : p ;
      p = a [ 18 ] & b [ 6 ] ? p + ( 60'h1 << 24 ) : p ;
      p = a [ 18 ] & b [ 7 ] ? p + ( 60'h1 << 25 ) : p ;
      p = a [ 18 ] & b [ 8 ] ? p + ( 60'h1 << 26 ) : p ;
      p = a [ 18 ] & b [ 9 ] ? p + ( 60'h1 << 27 ) : p ;
      p = a [ 18 ] & b [ 10 ] ? p + ( 60'h1 << 28 ) : p ;
      p = a [ 18 ] & b [ 11 ] ? p + ( 60'h1 << 29 ) : p ;
      p = a [ 18 ] & b [ 12 ] ? p + ( 60'h1 << 30 ) : p ;
      p = a [ 18 ] & b [ 13 ] ? p + ( 60'h1 << 31 ) : p ;
      p = a [ 18 ] & b [ 14 ] ? p + ( 60'h1 << 32 ) : p ;
      p = a [ 18 ] & b [ 15 ] ? p + ( 60'h1 << 33 ) : p ;
      p = a [ 18 ] & b [ 16 ] ? p + ( 60'h1 << 34 ) : p ;
      p = a [ 18 ] & b [ 17 ] ? p + ( 60'h1 << 35 ) : p ;
      p = a [ 18 ] & b [ 18 ] ? p + ( 60'h1 << 36 ) : p ;
      p = a [ 18 ] & b [ 19 ] ? p + ( 60'h1 << 37 ) : p ;
      p = a [ 18 ] & b [ 20 ] ? p + ( 60'h1 << 38 ) : p ;
      p = a [ 18 ] & b [ 21 ] ? p + ( 60'h1 << 39 ) : p ;
      p = a [ 18 ] & b [ 22 ] ? p + ( 60'h1 << 40 ) : p ;
      p = a [ 18 ] & b [ 23 ] ? p + ( 60'h1 << 41 ) : p ;
      p = a [ 18 ] & b [ 24 ] ? p + ( 60'h1 << 42 ) : p ;
      p = a [ 18 ] & b [ 25 ] ? p + ( 60'h1 << 43 ) : p ;
      p = a [ 18 ] & b [ 26 ] ? p + ( 60'h1 << 44 ) : p ;
      p = a [ 18 ] & b [ 27 ] ? p + ( 60'h1 << 45 ) : p ;
      p = a [ 18 ] & b [ 28 ] ? p + ( 60'h1 << 46 ) : p ;
      p = a [ 18 ] & b [ 29 ] ? p + ( 60'h1 << 47 ) : p ;
      p = a [ 18 ] & b [ 30 ] ? p + ( 60'h1 << 48 ) : p ;
      p = a [ 18 ] & b [ 31 ] ? p + ( 60'h1 << 49 ) : p ;
      p = a [ 18 ] & b [ 32 ] ? p + ( 60'h1 << 50 ) : p ;
      p = a [ 18 ] & b [ 33 ] ? p + ( 60'h1 << 51 ) : p ;
      p = a [ 18 ] & b [ 34 ] ? p + ( 60'h1 << 52 ) : p ;
      p = a [ 18 ] & b [ 35 ] ? p + ( 60'h1 << 53 ) : p ;
      p = a [ 18 ] & b [ 36 ] ? p + ( 60'h1 << 54 ) : p ;
      p = a [ 18 ] & b [ 37 ] ? p + ( 60'h1 << 55 ) : p ;
      p = a [ 18 ] & b [ 38 ] ? p + ( 60'h1 << 56 ) : p ;
      p = a [ 18 ] & b [ 39 ] ? p + ( 60'h1 << 57 ) : p ;
      p = a [ 18 ] & b [ 40 ] ? p + ( 60'h1 << 58 ) : p ;
      p = a [ 18 ] & b [ 41 ] ? p + ( 60'h1 << 59 ) : p ;

// Bit by Bit Multiply & Divide + Modulus
// Copyright © 2022 by Gregory Scott Callen
// All Rights Reserved.

      p = a [ 19 ] & b [ 0 ] ? p + ( 60'h1 << 19 ) : p ;
      p = a [ 19 ] & b [ 1 ] ? p + ( 60'h1 << 20 ) : p ;
      p = a [ 19 ] & b [ 2 ] ? p + ( 60'h1 << 21 ) : p ;
      p = a [ 19 ] & b [ 3 ] ? p + ( 60'h1 << 22 ) : p ;
      p = a [ 19 ] & b [ 4 ] ? p + ( 60'h1 << 23 ) : p ;
      p = a [ 19 ] & b [ 5 ] ? p + ( 60'h1 << 24 ) : p ;
      p = a [ 19 ] & b [ 6 ] ? p + ( 60'h1 << 25 ) : p ;
      p = a [ 19 ] & b [ 7 ] ? p + ( 60'h1 << 26 ) : p ;
      p = a [ 19 ] & b [ 8 ] ? p + ( 60'h1 << 27 ) : p ;
      p = a [ 19 ] & b [ 9 ] ? p + ( 60'h1 << 28 ) : p ;
      p = a [ 19 ] & b [ 10 ] ? p + ( 60'h1 << 29 ) : p ;
      p = a [ 19 ] & b [ 11 ] ? p + ( 60'h1 << 30 ) : p ;
      p = a [ 19 ] & b [ 12 ] ? p + ( 60'h1 << 31 ) : p ;
      p = a [ 19 ] & b [ 13 ] ? p + ( 60'h1 << 32 ) : p ;
      p = a [ 19 ] & b [ 14 ] ? p + ( 60'h1 << 33 ) : p ;
      p = a [ 19 ] & b [ 15 ] ? p + ( 60'h1 << 34 ) : p ;
      p = a [ 19 ] & b [ 16 ] ? p + ( 60'h1 << 35 ) : p ;
      p = a [ 19 ] & b [ 17 ] ? p + ( 60'h1 << 36 ) : p ;
      p = a [ 19 ] & b [ 18 ] ? p + ( 60'h1 << 37 ) : p ;
      p = a [ 19 ] & b [ 19 ] ? p + ( 60'h1 << 38 ) : p ;
      p = a [ 19 ] & b [ 20 ] ? p + ( 60'h1 << 39 ) : p ;
      p = a [ 19 ] & b [ 21 ] ? p + ( 60'h1 << 40 ) : p ;
      p = a [ 19 ] & b [ 22 ] ? p + ( 60'h1 << 41 ) : p ;
      p = a [ 19 ] & b [ 23 ] ? p + ( 60'h1 << 42 ) : p ;
      p = a [ 19 ] & b [ 24 ] ? p + ( 60'h1 << 43 ) : p ;
      p = a [ 19 ] & b [ 25 ] ? p + ( 60'h1 << 44 ) : p ;
      p = a [ 19 ] & b [ 26 ] ? p + ( 60'h1 << 45 ) : p ;
      p = a [ 19 ] & b [ 27 ] ? p + ( 60'h1 << 46 ) : p ;
      p = a [ 19 ] & b [ 28 ] ? p + ( 60'h1 << 47 ) : p ;
      p = a [ 19 ] & b [ 29 ] ? p + ( 60'h1 << 48 ) : p ;
      p = a [ 19 ] & b [ 30 ] ? p + ( 60'h1 << 49 ) : p ;
      p = a [ 19 ] & b [ 31 ] ? p + ( 60'h1 << 50 ) : p ;
      p = a [ 19 ] & b [ 32 ] ? p + ( 60'h1 << 51 ) : p ;
      p = a [ 19 ] & b [ 33 ] ? p + ( 60'h1 << 52 ) : p ;
      p = a [ 19 ] & b [ 34 ] ? p + ( 60'h1 << 53 ) : p ;
      p = a [ 19 ] & b [ 35 ] ? p + ( 60'h1 << 54 ) : p ;
      p = a [ 19 ] & b [ 36 ] ? p + ( 60'h1 << 55 ) : p ;
      p = a [ 19 ] & b [ 37 ] ? p + ( 60'h1 << 56 ) : p ;
      p = a [ 19 ] & b [ 38 ] ? p + ( 60'h1 << 57 ) : p ;
      p = a [ 19 ] & b [ 39 ] ? p + ( 60'h1 << 58 ) : p ;
      p = a [ 19 ] & b [ 40 ] ? p + ( 60'h1 << 59 ) : p ;

// Bit by Bit Multiply & Divide + Modulus
// Copyright © 2022 by Gregory Scott Callen
// All Rights Reserved.

      p = a [ 20 ] & b [ 0 ] ? p + ( 60'h1 << 20 ) : p ;
      p = a [ 20 ] & b [ 1 ] ? p + ( 60'h1 << 21 ) : p ;
      p = a [ 20 ] & b [ 2 ] ? p + ( 60'h1 << 22 ) : p ;
      p = a [ 20 ] & b [ 3 ] ? p + ( 60'h1 << 23 ) : p ;
      p = a [ 20 ] & b [ 4 ] ? p + ( 60'h1 << 24 ) : p ;
      p = a [ 20 ] & b [ 5 ] ? p + ( 60'h1 << 25 ) : p ;
      p = a [ 20 ] & b [ 6 ] ? p + ( 60'h1 << 26 ) : p ;
      p = a [ 20 ] & b [ 7 ] ? p + ( 60'h1 << 27 ) : p ;
      p = a [ 20 ] & b [ 8 ] ? p + ( 60'h1 << 28 ) : p ;
      p = a [ 20 ] & b [ 9 ] ? p + ( 60'h1 << 29 ) : p ;
      p = a [ 20 ] & b [ 10 ] ? p + ( 60'h1 << 30 ) : p ;
      p = a [ 20 ] & b [ 11 ] ? p + ( 60'h1 << 31 ) : p ;
      p = a [ 20 ] & b [ 12 ] ? p + ( 60'h1 << 32 ) : p ;
      p = a [ 20 ] & b [ 13 ] ? p + ( 60'h1 << 33 ) : p ;
      p = a [ 20 ] & b [ 14 ] ? p + ( 60'h1 << 34 ) : p ;
      p = a [ 20 ] & b [ 15 ] ? p + ( 60'h1 << 35 ) : p ;
      p = a [ 20 ] & b [ 16 ] ? p + ( 60'h1 << 36 ) : p ;
      p = a [ 20 ] & b [ 17 ] ? p + ( 60'h1 << 37 ) : p ;
      p = a [ 20 ] & b [ 18 ] ? p + ( 60'h1 << 38 ) : p ;
      p = a [ 20 ] & b [ 19 ] ? p + ( 60'h1 << 39 ) : p ;
      p = a [ 20 ] & b [ 20 ] ? p + ( 60'h1 << 40 ) : p ;
      p = a [ 20 ] & b [ 21 ] ? p + ( 60'h1 << 41 ) : p ;
      p = a [ 20 ] & b [ 22 ] ? p + ( 60'h1 << 42 ) : p ;
      p = a [ 20 ] & b [ 23 ] ? p + ( 60'h1 << 43 ) : p ;
      p = a [ 20 ] & b [ 24 ] ? p + ( 60'h1 << 44 ) : p ;
      p = a [ 20 ] & b [ 25 ] ? p + ( 60'h1 << 45 ) : p ;
      p = a [ 20 ] & b [ 26 ] ? p + ( 60'h1 << 46 ) : p ;
      p = a [ 20 ] & b [ 27 ] ? p + ( 60'h1 << 47 ) : p ;
      p = a [ 20 ] & b [ 28 ] ? p + ( 60'h1 << 48 ) : p ;
      p = a [ 20 ] & b [ 29 ] ? p + ( 60'h1 << 49 ) : p ;
      p = a [ 20 ] & b [ 30 ] ? p + ( 60'h1 << 50 ) : p ;
      p = a [ 20 ] & b [ 31 ] ? p + ( 60'h1 << 51 ) : p ;
      p = a [ 20 ] & b [ 32 ] ? p + ( 60'h1 << 52 ) : p ;
      p = a [ 20 ] & b [ 33 ] ? p + ( 60'h1 << 53 ) : p ;
      p = a [ 20 ] & b [ 34 ] ? p + ( 60'h1 << 54 ) : p ;
      p = a [ 20 ] & b [ 35 ] ? p + ( 60'h1 << 55 ) : p ;
      p = a [ 20 ] & b [ 36 ] ? p + ( 60'h1 << 56 ) : p ;
      p = a [ 20 ] & b [ 37 ] ? p + ( 60'h1 << 57 ) : p ;
      p = a [ 20 ] & b [ 38 ] ? p + ( 60'h1 << 58 ) : p ;
      p = a [ 20 ] & b [ 39 ] ? p + ( 60'h1 << 59 ) : p ;

// Bit by Bit Multiply & Divide + Modulus
// Copyright © 2022 by Gregory Scott Callen
// All Rights Reserved.

      p = a [ 21 ] & b [ 0 ] ? p + ( 60'h1 << 21 ) : p ;
      p = a [ 21 ] & b [ 1 ] ? p + ( 60'h1 << 22 ) : p ;
      p = a [ 21 ] & b [ 2 ] ? p + ( 60'h1 << 23 ) : p ;
      p = a [ 21 ] & b [ 3 ] ? p + ( 60'h1 << 24 ) : p ;
      p = a [ 21 ] & b [ 4 ] ? p + ( 60'h1 << 25 ) : p ;
      p = a [ 21 ] & b [ 5 ] ? p + ( 60'h1 << 26 ) : p ;
      p = a [ 21 ] & b [ 6 ] ? p + ( 60'h1 << 27 ) : p ;
      p = a [ 21 ] & b [ 7 ] ? p + ( 60'h1 << 28 ) : p ;
      p = a [ 21 ] & b [ 8 ] ? p + ( 60'h1 << 29 ) : p ;
      p = a [ 21 ] & b [ 9 ] ? p + ( 60'h1 << 30 ) : p ;
      p = a [ 21 ] & b [ 10 ] ? p + ( 60'h1 << 31 ) : p ;
      p = a [ 21 ] & b [ 11 ] ? p + ( 60'h1 << 32 ) : p ;
      p = a [ 21 ] & b [ 12 ] ? p + ( 60'h1 << 33 ) : p ;
      p = a [ 21 ] & b [ 13 ] ? p + ( 60'h1 << 34 ) : p ;
      p = a [ 21 ] & b [ 14 ] ? p + ( 60'h1 << 35 ) : p ;
      p = a [ 21 ] & b [ 15 ] ? p + ( 60'h1 << 36 ) : p ;
      p = a [ 21 ] & b [ 16 ] ? p + ( 60'h1 << 37 ) : p ;
      p = a [ 21 ] & b [ 17 ] ? p + ( 60'h1 << 38 ) : p ;
      p = a [ 21 ] & b [ 18 ] ? p + ( 60'h1 << 39 ) : p ;
      p = a [ 21 ] & b [ 19 ] ? p + ( 60'h1 << 40 ) : p ;
      p = a [ 21 ] & b [ 20 ] ? p + ( 60'h1 << 41 ) : p ;
      p = a [ 21 ] & b [ 21 ] ? p + ( 60'h1 << 42 ) : p ;
      p = a [ 21 ] & b [ 22 ] ? p + ( 60'h1 << 43 ) : p ;
      p = a [ 21 ] & b [ 23 ] ? p + ( 60'h1 << 44 ) : p ;
      p = a [ 21 ] & b [ 24 ] ? p + ( 60'h1 << 45 ) : p ;
      p = a [ 21 ] & b [ 25 ] ? p + ( 60'h1 << 46 ) : p ;
      p = a [ 21 ] & b [ 26 ] ? p + ( 60'h1 << 47 ) : p ;
      p = a [ 21 ] & b [ 27 ] ? p + ( 60'h1 << 48 ) : p ;
      p = a [ 21 ] & b [ 28 ] ? p + ( 60'h1 << 49 ) : p ;
      p = a [ 21 ] & b [ 29 ] ? p + ( 60'h1 << 50 ) : p ;
      p = a [ 21 ] & b [ 30 ] ? p + ( 60'h1 << 51 ) : p ;
      p = a [ 21 ] & b [ 31 ] ? p + ( 60'h1 << 52 ) : p ;
      p = a [ 21 ] & b [ 32 ] ? p + ( 60'h1 << 53 ) : p ;
      p = a [ 21 ] & b [ 33 ] ? p + ( 60'h1 << 54 ) : p ;
      p = a [ 21 ] & b [ 34 ] ? p + ( 60'h1 << 55 ) : p ;
      p = a [ 21 ] & b [ 35 ] ? p + ( 60'h1 << 56 ) : p ;
      p = a [ 21 ] & b [ 36 ] ? p + ( 60'h1 << 57 ) : p ;
      p = a [ 21 ] & b [ 37 ] ? p + ( 60'h1 << 58 ) : p ;
      p = a [ 21 ] & b [ 38 ] ? p + ( 60'h1 << 59 ) : p ;

// Bit by Bit Multiply & Divide + Modulus
// Copyright © 2022 by Gregory Scott Callen
// All Rights Reserved.

      p = a [ 22 ] & b [ 0 ] ? p + ( 60'h1 << 22 ) : p ;
      p = a [ 22 ] & b [ 1 ] ? p + ( 60'h1 << 23 ) : p ;
      p = a [ 22 ] & b [ 2 ] ? p + ( 60'h1 << 24 ) : p ;
      p = a [ 22 ] & b [ 3 ] ? p + ( 60'h1 << 25 ) : p ;
      p = a [ 22 ] & b [ 4 ] ? p + ( 60'h1 << 26 ) : p ;
      p = a [ 22 ] & b [ 5 ] ? p + ( 60'h1 << 27 ) : p ;
      p = a [ 22 ] & b [ 6 ] ? p + ( 60'h1 << 28 ) : p ;
      p = a [ 22 ] & b [ 7 ] ? p + ( 60'h1 << 29 ) : p ;
      p = a [ 22 ] & b [ 8 ] ? p + ( 60'h1 << 30 ) : p ;
      p = a [ 22 ] & b [ 9 ] ? p + ( 60'h1 << 31 ) : p ;
      p = a [ 22 ] & b [ 10 ] ? p + ( 60'h1 << 32 ) : p ;
      p = a [ 22 ] & b [ 11 ] ? p + ( 60'h1 << 33 ) : p ;
      p = a [ 22 ] & b [ 12 ] ? p + ( 60'h1 << 34 ) : p ;
      p = a [ 22 ] & b [ 13 ] ? p + ( 60'h1 << 35 ) : p ;
      p = a [ 22 ] & b [ 14 ] ? p + ( 60'h1 << 36 ) : p ;
      p = a [ 22 ] & b [ 15 ] ? p + ( 60'h1 << 37 ) : p ;
      p = a [ 22 ] & b [ 16 ] ? p + ( 60'h1 << 38 ) : p ;
      p = a [ 22 ] & b [ 17 ] ? p + ( 60'h1 << 39 ) : p ;
      p = a [ 22 ] & b [ 18 ] ? p + ( 60'h1 << 40 ) : p ;
      p = a [ 22 ] & b [ 19 ] ? p + ( 60'h1 << 41 ) : p ;
      p = a [ 22 ] & b [ 20 ] ? p + ( 60'h1 << 42 ) : p ;
      p = a [ 22 ] & b [ 21 ] ? p + ( 60'h1 << 43 ) : p ;
      p = a [ 22 ] & b [ 22 ] ? p + ( 60'h1 << 44 ) : p ;
      p = a [ 22 ] & b [ 23 ] ? p + ( 60'h1 << 45 ) : p ;
      p = a [ 22 ] & b [ 24 ] ? p + ( 60'h1 << 46 ) : p ;
      p = a [ 22 ] & b [ 25 ] ? p + ( 60'h1 << 47 ) : p ;
      p = a [ 22 ] & b [ 26 ] ? p + ( 60'h1 << 48 ) : p ;
      p = a [ 22 ] & b [ 27 ] ? p + ( 60'h1 << 49 ) : p ;
      p = a [ 22 ] & b [ 28 ] ? p + ( 60'h1 << 50 ) : p ;
      p = a [ 22 ] & b [ 29 ] ? p + ( 60'h1 << 51 ) : p ;
      p = a [ 22 ] & b [ 30 ] ? p + ( 60'h1 << 52 ) : p ;
      p = a [ 22 ] & b [ 31 ] ? p + ( 60'h1 << 53 ) : p ;
      p = a [ 22 ] & b [ 32 ] ? p + ( 60'h1 << 54 ) : p ;
      p = a [ 22 ] & b [ 33 ] ? p + ( 60'h1 << 55 ) : p ;
      p = a [ 22 ] & b [ 34 ] ? p + ( 60'h1 << 56 ) : p ;
      p = a [ 22 ] & b [ 35 ] ? p + ( 60'h1 << 57 ) : p ;
      p = a [ 22 ] & b [ 36 ] ? p + ( 60'h1 << 58 ) : p ;
      p = a [ 22 ] & b [ 37 ] ? p + ( 60'h1 << 59 ) : p ;

// Bit by Bit Multiply & Divide + Modulus
// Copyright © 2022 by Gregory Scott Callen
// All Rights Reserved.

      p = a [ 23 ] & b [ 0 ] ? p + ( 60'h1 << 23 ) : p ;
      p = a [ 23 ] & b [ 1 ] ? p + ( 60'h1 << 24 ) : p ;
      p = a [ 23 ] & b [ 2 ] ? p + ( 60'h1 << 25 ) : p ;
      p = a [ 23 ] & b [ 3 ] ? p + ( 60'h1 << 26 ) : p ;
      p = a [ 23 ] & b [ 4 ] ? p + ( 60'h1 << 27 ) : p ;
      p = a [ 23 ] & b [ 5 ] ? p + ( 60'h1 << 28 ) : p ;
      p = a [ 23 ] & b [ 6 ] ? p + ( 60'h1 << 29 ) : p ;
      p = a [ 23 ] & b [ 7 ] ? p + ( 60'h1 << 30 ) : p ;
      p = a [ 23 ] & b [ 8 ] ? p + ( 60'h1 << 31 ) : p ;
      p = a [ 23 ] & b [ 9 ] ? p + ( 60'h1 << 32 ) : p ;
      p = a [ 23 ] & b [ 10 ] ? p + ( 60'h1 << 33 ) : p ;
      p = a [ 23 ] & b [ 11 ] ? p + ( 60'h1 << 34 ) : p ;
      p = a [ 23 ] & b [ 12 ] ? p + ( 60'h1 << 35 ) : p ;
      p = a [ 23 ] & b [ 13 ] ? p + ( 60'h1 << 36 ) : p ;
      p = a [ 23 ] & b [ 14 ] ? p + ( 60'h1 << 37 ) : p ;
      p = a [ 23 ] & b [ 15 ] ? p + ( 60'h1 << 38 ) : p ;
      p = a [ 23 ] & b [ 16 ] ? p + ( 60'h1 << 39 ) : p ;
      p = a [ 23 ] & b [ 17 ] ? p + ( 60'h1 << 40 ) : p ;
      p = a [ 23 ] & b [ 18 ] ? p + ( 60'h1 << 41 ) : p ;
      p = a [ 23 ] & b [ 19 ] ? p + ( 60'h1 << 42 ) : p ;
      p = a [ 23 ] & b [ 20 ] ? p + ( 60'h1 << 43 ) : p ;
      p = a [ 23 ] & b [ 21 ] ? p + ( 60'h1 << 44 ) : p ;
      p = a [ 23 ] & b [ 22 ] ? p + ( 60'h1 << 45 ) : p ;
      p = a [ 23 ] & b [ 23 ] ? p + ( 60'h1 << 46 ) : p ;
      p = a [ 23 ] & b [ 24 ] ? p + ( 60'h1 << 47 ) : p ;
      p = a [ 23 ] & b [ 25 ] ? p + ( 60'h1 << 48 ) : p ;
      p = a [ 23 ] & b [ 26 ] ? p + ( 60'h1 << 49 ) : p ;
      p = a [ 23 ] & b [ 27 ] ? p + ( 60'h1 << 50 ) : p ;
      p = a [ 23 ] & b [ 28 ] ? p + ( 60'h1 << 51 ) : p ;
      p = a [ 23 ] & b [ 29 ] ? p + ( 60'h1 << 52 ) : p ;
      p = a [ 23 ] & b [ 30 ] ? p + ( 60'h1 << 53 ) : p ;
      p = a [ 23 ] & b [ 31 ] ? p + ( 60'h1 << 54 ) : p ;
      p = a [ 23 ] & b [ 32 ] ? p + ( 60'h1 << 55 ) : p ;
      p = a [ 23 ] & b [ 33 ] ? p + ( 60'h1 << 56 ) : p ;
      p = a [ 23 ] & b [ 34 ] ? p + ( 60'h1 << 57 ) : p ;
      p = a [ 23 ] & b [ 35 ] ? p + ( 60'h1 << 58 ) : p ;
      p = a [ 23 ] & b [ 36 ] ? p + ( 60'h1 << 59 ) : p ;

// Bit by Bit Multiply & Divide + Modulus
// Copyright © 2022 by Gregory Scott Callen
// All Rights Reserved.

      p = a [ 24 ] & b [ 0 ] ? p + ( 60'h1 << 24 ) : p ;
      p = a [ 24 ] & b [ 1 ] ? p + ( 60'h1 << 25 ) : p ;
      p = a [ 24 ] & b [ 2 ] ? p + ( 60'h1 << 26 ) : p ;
      p = a [ 24 ] & b [ 3 ] ? p + ( 60'h1 << 27 ) : p ;
      p = a [ 24 ] & b [ 4 ] ? p + ( 60'h1 << 28 ) : p ;
      p = a [ 24 ] & b [ 5 ] ? p + ( 60'h1 << 29 ) : p ;
      p = a [ 24 ] & b [ 6 ] ? p + ( 60'h1 << 30 ) : p ;
      p = a [ 24 ] & b [ 7 ] ? p + ( 60'h1 << 31 ) : p ;
      p = a [ 24 ] & b [ 8 ] ? p + ( 60'h1 << 32 ) : p ;
      p = a [ 24 ] & b [ 9 ] ? p + ( 60'h1 << 33 ) : p ;
      p = a [ 24 ] & b [ 10 ] ? p + ( 60'h1 << 34 ) : p ;
      p = a [ 24 ] & b [ 11 ] ? p + ( 60'h1 << 35 ) : p ;
      p = a [ 24 ] & b [ 12 ] ? p + ( 60'h1 << 36 ) : p ;
      p = a [ 24 ] & b [ 13 ] ? p + ( 60'h1 << 37 ) : p ;
      p = a [ 24 ] & b [ 14 ] ? p + ( 60'h1 << 38 ) : p ;
      p = a [ 24 ] & b [ 15 ] ? p + ( 60'h1 << 39 ) : p ;
      p = a [ 24 ] & b [ 16 ] ? p + ( 60'h1 << 40 ) : p ;
      p = a [ 24 ] & b [ 17 ] ? p + ( 60'h1 << 41 ) : p ;
      p = a [ 24 ] & b [ 18 ] ? p + ( 60'h1 << 42 ) : p ;
      p = a [ 24 ] & b [ 19 ] ? p + ( 60'h1 << 43 ) : p ;
      p = a [ 24 ] & b [ 20 ] ? p + ( 60'h1 << 44 ) : p ;
      p = a [ 24 ] & b [ 21 ] ? p + ( 60'h1 << 45 ) : p ;
      p = a [ 24 ] & b [ 22 ] ? p + ( 60'h1 << 46 ) : p ;
      p = a [ 24 ] & b [ 23 ] ? p + ( 60'h1 << 47 ) : p ;
      p = a [ 24 ] & b [ 24 ] ? p + ( 60'h1 << 48 ) : p ;
      p = a [ 24 ] & b [ 25 ] ? p + ( 60'h1 << 49 ) : p ;
      p = a [ 24 ] & b [ 26 ] ? p + ( 60'h1 << 50 ) : p ;
      p = a [ 24 ] & b [ 27 ] ? p + ( 60'h1 << 51 ) : p ;
      p = a [ 24 ] & b [ 28 ] ? p + ( 60'h1 << 52 ) : p ;
      p = a [ 24 ] & b [ 29 ] ? p + ( 60'h1 << 53 ) : p ;
      p = a [ 24 ] & b [ 30 ] ? p + ( 60'h1 << 54 ) : p ;
      p = a [ 24 ] & b [ 31 ] ? p + ( 60'h1 << 55 ) : p ;
      p = a [ 24 ] & b [ 32 ] ? p + ( 60'h1 << 56 ) : p ;
      p = a [ 24 ] & b [ 33 ] ? p + ( 60'h1 << 57 ) : p ;
      p = a [ 24 ] & b [ 34 ] ? p + ( 60'h1 << 58 ) : p ;
      p = a [ 24 ] & b [ 35 ] ? p + ( 60'h1 << 59 ) : p ;

// Bit by Bit Multiply & Divide + Modulus
// Copyright © 2022 by Gregory Scott Callen
// All Rights Reserved.

      p = a [ 25 ] & b [ 0 ] ? p + ( 60'h1 << 25 ) : p ;
      p = a [ 25 ] & b [ 1 ] ? p + ( 60'h1 << 26 ) : p ;
      p = a [ 25 ] & b [ 2 ] ? p + ( 60'h1 << 27 ) : p ;
      p = a [ 25 ] & b [ 3 ] ? p + ( 60'h1 << 28 ) : p ;
      p = a [ 25 ] & b [ 4 ] ? p + ( 60'h1 << 29 ) : p ;
      p = a [ 25 ] & b [ 5 ] ? p + ( 60'h1 << 30 ) : p ;
      p = a [ 25 ] & b [ 6 ] ? p + ( 60'h1 << 31 ) : p ;
      p = a [ 25 ] & b [ 7 ] ? p + ( 60'h1 << 32 ) : p ;
      p = a [ 25 ] & b [ 8 ] ? p + ( 60'h1 << 33 ) : p ;
      p = a [ 25 ] & b [ 9 ] ? p + ( 60'h1 << 34 ) : p ;
      p = a [ 25 ] & b [ 10 ] ? p + ( 60'h1 << 35 ) : p ;
      p = a [ 25 ] & b [ 11 ] ? p + ( 60'h1 << 36 ) : p ;
      p = a [ 25 ] & b [ 12 ] ? p + ( 60'h1 << 37 ) : p ;
      p = a [ 25 ] & b [ 13 ] ? p + ( 60'h1 << 38 ) : p ;
      p = a [ 25 ] & b [ 14 ] ? p + ( 60'h1 << 39 ) : p ;
      p = a [ 25 ] & b [ 15 ] ? p + ( 60'h1 << 40 ) : p ;
      p = a [ 25 ] & b [ 16 ] ? p + ( 60'h1 << 41 ) : p ;
      p = a [ 25 ] & b [ 17 ] ? p + ( 60'h1 << 42 ) : p ;
      p = a [ 25 ] & b [ 18 ] ? p + ( 60'h1 << 43 ) : p ;
      p = a [ 25 ] & b [ 19 ] ? p + ( 60'h1 << 44 ) : p ;
      p = a [ 25 ] & b [ 20 ] ? p + ( 60'h1 << 45 ) : p ;
      p = a [ 25 ] & b [ 21 ] ? p + ( 60'h1 << 46 ) : p ;
      p = a [ 25 ] & b [ 22 ] ? p + ( 60'h1 << 47 ) : p ;
      p = a [ 25 ] & b [ 23 ] ? p + ( 60'h1 << 48 ) : p ;
      p = a [ 25 ] & b [ 24 ] ? p + ( 60'h1 << 49 ) : p ;
      p = a [ 25 ] & b [ 25 ] ? p + ( 60'h1 << 50 ) : p ;
      p = a [ 25 ] & b [ 26 ] ? p + ( 60'h1 << 51 ) : p ;
      p = a [ 25 ] & b [ 27 ] ? p + ( 60'h1 << 52 ) : p ;
      p = a [ 25 ] & b [ 28 ] ? p + ( 60'h1 << 53 ) : p ;
      p = a [ 25 ] & b [ 29 ] ? p + ( 60'h1 << 54 ) : p ;
      p = a [ 25 ] & b [ 30 ] ? p + ( 60'h1 << 55 ) : p ;
      p = a [ 25 ] & b [ 31 ] ? p + ( 60'h1 << 56 ) : p ;
      p = a [ 25 ] & b [ 32 ] ? p + ( 60'h1 << 57 ) : p ;
      p = a [ 25 ] & b [ 33 ] ? p + ( 60'h1 << 58 ) : p ;
      p = a [ 25 ] & b [ 34 ] ? p + ( 60'h1 << 59 ) : p ;

// Bit by Bit Multiply & Divide + Modulus
// Copyright © 2022 by Gregory Scott Callen
// All Rights Reserved.

      p = a [ 26 ] & b [ 0 ] ? p + ( 60'h1 << 26 ) : p ;
      p = a [ 26 ] & b [ 1 ] ? p + ( 60'h1 << 27 ) : p ;
      p = a [ 26 ] & b [ 2 ] ? p + ( 60'h1 << 28 ) : p ;
      p = a [ 26 ] & b [ 3 ] ? p + ( 60'h1 << 29 ) : p ;
      p = a [ 26 ] & b [ 4 ] ? p + ( 60'h1 << 30 ) : p ;
      p = a [ 26 ] & b [ 5 ] ? p + ( 60'h1 << 31 ) : p ;
      p = a [ 26 ] & b [ 6 ] ? p + ( 60'h1 << 32 ) : p ;
      p = a [ 26 ] & b [ 7 ] ? p + ( 60'h1 << 33 ) : p ;
      p = a [ 26 ] & b [ 8 ] ? p + ( 60'h1 << 34 ) : p ;
      p = a [ 26 ] & b [ 9 ] ? p + ( 60'h1 << 35 ) : p ;
      p = a [ 26 ] & b [ 10 ] ? p + ( 60'h1 << 36 ) : p ;
      p = a [ 26 ] & b [ 11 ] ? p + ( 60'h1 << 37 ) : p ;
      p = a [ 26 ] & b [ 12 ] ? p + ( 60'h1 << 38 ) : p ;
      p = a [ 26 ] & b [ 13 ] ? p + ( 60'h1 << 39 ) : p ;
      p = a [ 26 ] & b [ 14 ] ? p + ( 60'h1 << 40 ) : p ;
      p = a [ 26 ] & b [ 15 ] ? p + ( 60'h1 << 41 ) : p ;
      p = a [ 26 ] & b [ 16 ] ? p + ( 60'h1 << 42 ) : p ;
      p = a [ 26 ] & b [ 17 ] ? p + ( 60'h1 << 43 ) : p ;
      p = a [ 26 ] & b [ 18 ] ? p + ( 60'h1 << 44 ) : p ;
      p = a [ 26 ] & b [ 19 ] ? p + ( 60'h1 << 45 ) : p ;
      p = a [ 26 ] & b [ 20 ] ? p + ( 60'h1 << 46 ) : p ;
      p = a [ 26 ] & b [ 21 ] ? p + ( 60'h1 << 47 ) : p ;
      p = a [ 26 ] & b [ 22 ] ? p + ( 60'h1 << 48 ) : p ;
      p = a [ 26 ] & b [ 23 ] ? p + ( 60'h1 << 49 ) : p ;
      p = a [ 26 ] & b [ 24 ] ? p + ( 60'h1 << 50 ) : p ;
      p = a [ 26 ] & b [ 25 ] ? p + ( 60'h1 << 51 ) : p ;
      p = a [ 26 ] & b [ 26 ] ? p + ( 60'h1 << 52 ) : p ;
      p = a [ 26 ] & b [ 27 ] ? p + ( 60'h1 << 53 ) : p ;
      p = a [ 26 ] & b [ 28 ] ? p + ( 60'h1 << 54 ) : p ;
      p = a [ 26 ] & b [ 29 ] ? p + ( 60'h1 << 55 ) : p ;
      p = a [ 26 ] & b [ 30 ] ? p + ( 60'h1 << 56 ) : p ;
      p = a [ 26 ] & b [ 31 ] ? p + ( 60'h1 << 57 ) : p ;
      p = a [ 26 ] & b [ 32 ] ? p + ( 60'h1 << 58 ) : p ;
      p = a [ 26 ] & b [ 33 ] ? p + ( 60'h1 << 59 ) : p ;

// Bit by Bit Multiply & Divide + Modulus
// Copyright © 2022 by Gregory Scott Callen
// All Rights Reserved.

      p = a [ 27 ] & b [ 0 ] ? p + ( 60'h1 << 27 ) : p ;
      p = a [ 27 ] & b [ 1 ] ? p + ( 60'h1 << 28 ) : p ;
      p = a [ 27 ] & b [ 2 ] ? p + ( 60'h1 << 29 ) : p ;
      p = a [ 27 ] & b [ 3 ] ? p + ( 60'h1 << 30 ) : p ;
      p = a [ 27 ] & b [ 4 ] ? p + ( 60'h1 << 31 ) : p ;
      p = a [ 27 ] & b [ 5 ] ? p + ( 60'h1 << 32 ) : p ;
      p = a [ 27 ] & b [ 6 ] ? p + ( 60'h1 << 33 ) : p ;
      p = a [ 27 ] & b [ 7 ] ? p + ( 60'h1 << 34 ) : p ;
      p = a [ 27 ] & b [ 8 ] ? p + ( 60'h1 << 35 ) : p ;
      p = a [ 27 ] & b [ 9 ] ? p + ( 60'h1 << 36 ) : p ;
      p = a [ 27 ] & b [ 10 ] ? p + ( 60'h1 << 37 ) : p ;
      p = a [ 27 ] & b [ 11 ] ? p + ( 60'h1 << 38 ) : p ;
      p = a [ 27 ] & b [ 12 ] ? p + ( 60'h1 << 39 ) : p ;
      p = a [ 27 ] & b [ 13 ] ? p + ( 60'h1 << 40 ) : p ;
      p = a [ 27 ] & b [ 14 ] ? p + ( 60'h1 << 41 ) : p ;
      p = a [ 27 ] & b [ 15 ] ? p + ( 60'h1 << 42 ) : p ;
      p = a [ 27 ] & b [ 16 ] ? p + ( 60'h1 << 43 ) : p ;
      p = a [ 27 ] & b [ 17 ] ? p + ( 60'h1 << 44 ) : p ;
      p = a [ 27 ] & b [ 18 ] ? p + ( 60'h1 << 45 ) : p ;
      p = a [ 27 ] & b [ 19 ] ? p + ( 60'h1 << 46 ) : p ;
      p = a [ 27 ] & b [ 20 ] ? p + ( 60'h1 << 47 ) : p ;
      p = a [ 27 ] & b [ 21 ] ? p + ( 60'h1 << 48 ) : p ;
      p = a [ 27 ] & b [ 22 ] ? p + ( 60'h1 << 49 ) : p ;
      p = a [ 27 ] & b [ 23 ] ? p + ( 60'h1 << 50 ) : p ;
      p = a [ 27 ] & b [ 24 ] ? p + ( 60'h1 << 51 ) : p ;
      p = a [ 27 ] & b [ 25 ] ? p + ( 60'h1 << 52 ) : p ;
      p = a [ 27 ] & b [ 26 ] ? p + ( 60'h1 << 53 ) : p ;
      p = a [ 27 ] & b [ 27 ] ? p + ( 60'h1 << 54 ) : p ;
      p = a [ 27 ] & b [ 28 ] ? p + ( 60'h1 << 55 ) : p ;
      p = a [ 27 ] & b [ 29 ] ? p + ( 60'h1 << 56 ) : p ;
      p = a [ 27 ] & b [ 30 ] ? p + ( 60'h1 << 57 ) : p ;
      p = a [ 27 ] & b [ 31 ] ? p + ( 60'h1 << 58 ) : p ;
      p = a [ 27 ] & b [ 32 ] ? p + ( 60'h1 << 59 ) : p ;

// Bit by Bit Multiply & Divide + Modulus
// Copyright © 2022 by Gregory Scott Callen
// All Rights Reserved.

      p = a [ 28 ] & b [ 0 ] ? p + ( 60'h1 << 28 ) : p ;
      p = a [ 28 ] & b [ 1 ] ? p + ( 60'h1 << 29 ) : p ;
      p = a [ 28 ] & b [ 2 ] ? p + ( 60'h1 << 30 ) : p ;
      p = a [ 28 ] & b [ 3 ] ? p + ( 60'h1 << 31 ) : p ;
      p = a [ 28 ] & b [ 4 ] ? p + ( 60'h1 << 32 ) : p ;
      p = a [ 28 ] & b [ 5 ] ? p + ( 60'h1 << 33 ) : p ;
      p = a [ 28 ] & b [ 6 ] ? p + ( 60'h1 << 34 ) : p ;
      p = a [ 28 ] & b [ 7 ] ? p + ( 60'h1 << 35 ) : p ;
      p = a [ 28 ] & b [ 8 ] ? p + ( 60'h1 << 36 ) : p ;
      p = a [ 28 ] & b [ 9 ] ? p + ( 60'h1 << 37 ) : p ;
      p = a [ 28 ] & b [ 10 ] ? p + ( 60'h1 << 38 ) : p ;
      p = a [ 28 ] & b [ 11 ] ? p + ( 60'h1 << 39 ) : p ;
      p = a [ 28 ] & b [ 12 ] ? p + ( 60'h1 << 40 ) : p ;
      p = a [ 28 ] & b [ 13 ] ? p + ( 60'h1 << 41 ) : p ;
      p = a [ 28 ] & b [ 14 ] ? p + ( 60'h1 << 42 ) : p ;
      p = a [ 28 ] & b [ 15 ] ? p + ( 60'h1 << 43 ) : p ;
      p = a [ 28 ] & b [ 16 ] ? p + ( 60'h1 << 44 ) : p ;
      p = a [ 28 ] & b [ 17 ] ? p + ( 60'h1 << 45 ) : p ;
      p = a [ 28 ] & b [ 18 ] ? p + ( 60'h1 << 46 ) : p ;
      p = a [ 28 ] & b [ 19 ] ? p + ( 60'h1 << 47 ) : p ;
      p = a [ 28 ] & b [ 20 ] ? p + ( 60'h1 << 48 ) : p ;
      p = a [ 28 ] & b [ 21 ] ? p + ( 60'h1 << 49 ) : p ;
      p = a [ 28 ] & b [ 22 ] ? p + ( 60'h1 << 50 ) : p ;
      p = a [ 28 ] & b [ 23 ] ? p + ( 60'h1 << 51 ) : p ;
      p = a [ 28 ] & b [ 24 ] ? p + ( 60'h1 << 52 ) : p ;
      p = a [ 28 ] & b [ 25 ] ? p + ( 60'h1 << 53 ) : p ;
      p = a [ 28 ] & b [ 26 ] ? p + ( 60'h1 << 54 ) : p ;
      p = a [ 28 ] & b [ 27 ] ? p + ( 60'h1 << 55 ) : p ;
      p = a [ 28 ] & b [ 28 ] ? p + ( 60'h1 << 56 ) : p ;
      p = a [ 28 ] & b [ 29 ] ? p + ( 60'h1 << 57 ) : p ;
      p = a [ 28 ] & b [ 30 ] ? p + ( 60'h1 << 58 ) : p ;
      p = a [ 28 ] & b [ 31 ] ? p + ( 60'h1 << 59 ) : p ;

// Bit by Bit Multiply & Divide + Modulus
// Copyright © 2022 by Gregory Scott Callen
// All Rights Reserved.

      p = a [ 29 ] & b [ 0 ] ? p + ( 60'h1 << 29 ) : p ;
      p = a [ 29 ] & b [ 1 ] ? p + ( 60'h1 << 30 ) : p ;
      p = a [ 29 ] & b [ 2 ] ? p + ( 60'h1 << 31 ) : p ;
      p = a [ 29 ] & b [ 3 ] ? p + ( 60'h1 << 32 ) : p ;
      p = a [ 29 ] & b [ 4 ] ? p + ( 60'h1 << 33 ) : p ;
      p = a [ 29 ] & b [ 5 ] ? p + ( 60'h1 << 34 ) : p ;
      p = a [ 29 ] & b [ 6 ] ? p + ( 60'h1 << 35 ) : p ;
      p = a [ 29 ] & b [ 7 ] ? p + ( 60'h1 << 36 ) : p ;
      p = a [ 29 ] & b [ 8 ] ? p + ( 60'h1 << 37 ) : p ;
      p = a [ 29 ] & b [ 9 ] ? p + ( 60'h1 << 38 ) : p ;
      p = a [ 29 ] & b [ 10 ] ? p + ( 60'h1 << 39 ) : p ;
      p = a [ 29 ] & b [ 11 ] ? p + ( 60'h1 << 40 ) : p ;
      p = a [ 29 ] & b [ 12 ] ? p + ( 60'h1 << 41 ) : p ;
      p = a [ 29 ] & b [ 13 ] ? p + ( 60'h1 << 42 ) : p ;
      p = a [ 29 ] & b [ 14 ] ? p + ( 60'h1 << 43 ) : p ;
      p = a [ 29 ] & b [ 15 ] ? p + ( 60'h1 << 44 ) : p ;
      p = a [ 29 ] & b [ 16 ] ? p + ( 60'h1 << 45 ) : p ;
      p = a [ 29 ] & b [ 17 ] ? p + ( 60'h1 << 46 ) : p ;
      p = a [ 29 ] & b [ 18 ] ? p + ( 60'h1 << 47 ) : p ;
      p = a [ 29 ] & b [ 19 ] ? p + ( 60'h1 << 48 ) : p ;
      p = a [ 29 ] & b [ 20 ] ? p + ( 60'h1 << 49 ) : p ;
      p = a [ 29 ] & b [ 21 ] ? p + ( 60'h1 << 50 ) : p ;
      p = a [ 29 ] & b [ 22 ] ? p + ( 60'h1 << 51 ) : p ;
      p = a [ 29 ] & b [ 23 ] ? p + ( 60'h1 << 52 ) : p ;
      p = a [ 29 ] & b [ 24 ] ? p + ( 60'h1 << 53 ) : p ;
      p = a [ 29 ] & b [ 25 ] ? p + ( 60'h1 << 54 ) : p ;
      p = a [ 29 ] & b [ 26 ] ? p + ( 60'h1 << 55 ) : p ;
      p = a [ 29 ] & b [ 27 ] ? p + ( 60'h1 << 56 ) : p ;
      p = a [ 29 ] & b [ 28 ] ? p + ( 60'h1 << 57 ) : p ;
      p = a [ 29 ] & b [ 29 ] ? p + ( 60'h1 << 58 ) : p ;
      p = a [ 29 ] & b [ 30 ] ? p + ( 60'h1 << 59 ) : p ;

// Bit by Bit Multiply & Divide + Modulus
// Copyright © 2022 by Gregory Scott Callen
// All Rights Reserved.

      p = a [ 30 ] & b [ 0 ] ? p + ( 60'h1 << 30 ) : p ;
      p = a [ 30 ] & b [ 1 ] ? p + ( 60'h1 << 31 ) : p ;
      p = a [ 30 ] & b [ 2 ] ? p + ( 60'h1 << 32 ) : p ;
      p = a [ 30 ] & b [ 3 ] ? p + ( 60'h1 << 33 ) : p ;
      p = a [ 30 ] & b [ 4 ] ? p + ( 60'h1 << 34 ) : p ;
      p = a [ 30 ] & b [ 5 ] ? p + ( 60'h1 << 35 ) : p ;
      p = a [ 30 ] & b [ 6 ] ? p + ( 60'h1 << 36 ) : p ;
      p = a [ 30 ] & b [ 7 ] ? p + ( 60'h1 << 37 ) : p ;
      p = a [ 30 ] & b [ 8 ] ? p + ( 60'h1 << 38 ) : p ;
      p = a [ 30 ] & b [ 9 ] ? p + ( 60'h1 << 39 ) : p ;
      p = a [ 30 ] & b [ 10 ] ? p + ( 60'h1 << 40 ) : p ;
      p = a [ 30 ] & b [ 11 ] ? p + ( 60'h1 << 41 ) : p ;
      p = a [ 30 ] & b [ 12 ] ? p + ( 60'h1 << 42 ) : p ;
      p = a [ 30 ] & b [ 13 ] ? p + ( 60'h1 << 43 ) : p ;
      p = a [ 30 ] & b [ 14 ] ? p + ( 60'h1 << 44 ) : p ;
      p = a [ 30 ] & b [ 15 ] ? p + ( 60'h1 << 45 ) : p ;
      p = a [ 30 ] & b [ 16 ] ? p + ( 60'h1 << 46 ) : p ;
      p = a [ 30 ] & b [ 17 ] ? p + ( 60'h1 << 47 ) : p ;
      p = a [ 30 ] & b [ 18 ] ? p + ( 60'h1 << 48 ) : p ;
      p = a [ 30 ] & b [ 19 ] ? p + ( 60'h1 << 49 ) : p ;
      p = a [ 30 ] & b [ 20 ] ? p + ( 60'h1 << 50 ) : p ;
      p = a [ 30 ] & b [ 21 ] ? p + ( 60'h1 << 51 ) : p ;
      p = a [ 30 ] & b [ 22 ] ? p + ( 60'h1 << 52 ) : p ;
      p = a [ 30 ] & b [ 23 ] ? p + ( 60'h1 << 53 ) : p ;
      p = a [ 30 ] & b [ 24 ] ? p + ( 60'h1 << 54 ) : p ;
      p = a [ 30 ] & b [ 25 ] ? p + ( 60'h1 << 55 ) : p ;
      p = a [ 30 ] & b [ 26 ] ? p + ( 60'h1 << 56 ) : p ;
      p = a [ 30 ] & b [ 27 ] ? p + ( 60'h1 << 57 ) : p ;
      p = a [ 30 ] & b [ 28 ] ? p + ( 60'h1 << 58 ) : p ;
      p = a [ 30 ] & b [ 29 ] ? p + ( 60'h1 << 59 ) : p ;

// Bit by Bit Multiply & Divide + Modulus
// Copyright © 2022 by Gregory Scott Callen
// All Rights Reserved.

      p = a [ 31 ] & b [ 0 ] ? p + ( 60'h1 << 31 ) : p ;
      p = a [ 31 ] & b [ 1 ] ? p + ( 60'h1 << 32 ) : p ;
      p = a [ 31 ] & b [ 2 ] ? p + ( 60'h1 << 33 ) : p ;
      p = a [ 31 ] & b [ 3 ] ? p + ( 60'h1 << 34 ) : p ;
      p = a [ 31 ] & b [ 4 ] ? p + ( 60'h1 << 35 ) : p ;
      p = a [ 31 ] & b [ 5 ] ? p + ( 60'h1 << 36 ) : p ;
      p = a [ 31 ] & b [ 6 ] ? p + ( 60'h1 << 37 ) : p ;
      p = a [ 31 ] & b [ 7 ] ? p + ( 60'h1 << 38 ) : p ;
      p = a [ 31 ] & b [ 8 ] ? p + ( 60'h1 << 39 ) : p ;
      p = a [ 31 ] & b [ 9 ] ? p + ( 60'h1 << 40 ) : p ;
      p = a [ 31 ] & b [ 10 ] ? p + ( 60'h1 << 41 ) : p ;
      p = a [ 31 ] & b [ 11 ] ? p + ( 60'h1 << 42 ) : p ;
      p = a [ 31 ] & b [ 12 ] ? p + ( 60'h1 << 43 ) : p ;
      p = a [ 31 ] & b [ 13 ] ? p + ( 60'h1 << 44 ) : p ;
      p = a [ 31 ] & b [ 14 ] ? p + ( 60'h1 << 45 ) : p ;
      p = a [ 31 ] & b [ 15 ] ? p + ( 60'h1 << 46 ) : p ;
      p = a [ 31 ] & b [ 16 ] ? p + ( 60'h1 << 47 ) : p ;
      p = a [ 31 ] & b [ 17 ] ? p + ( 60'h1 << 48 ) : p ;
      p = a [ 31 ] & b [ 18 ] ? p + ( 60'h1 << 49 ) : p ;
      p = a [ 31 ] & b [ 19 ] ? p + ( 60'h1 << 50 ) : p ;
      p = a [ 31 ] & b [ 20 ] ? p + ( 60'h1 << 51 ) : p ;
      p = a [ 31 ] & b [ 21 ] ? p + ( 60'h1 << 52 ) : p ;
      p = a [ 31 ] & b [ 22 ] ? p + ( 60'h1 << 53 ) : p ;
      p = a [ 31 ] & b [ 23 ] ? p + ( 60'h1 << 54 ) : p ;
      p = a [ 31 ] & b [ 24 ] ? p + ( 60'h1 << 55 ) : p ;
      p = a [ 31 ] & b [ 25 ] ? p + ( 60'h1 << 56 ) : p ;
      p = a [ 31 ] & b [ 26 ] ? p + ( 60'h1 << 57 ) : p ;
      p = a [ 31 ] & b [ 27 ] ? p + ( 60'h1 << 58 ) : p ;
      p = a [ 31 ] & b [ 28 ] ? p + ( 60'h1 << 59 ) : p ;

// Bit by Bit Multiply & Divide + Modulus
// Copyright © 2022 by Gregory Scott Callen
// All Rights Reserved.

      p = a [ 32 ] & b [ 0 ] ? p + ( 60'h1 << 32 ) : p ;
      p = a [ 32 ] & b [ 1 ] ? p + ( 60'h1 << 33 ) : p ;
      p = a [ 32 ] & b [ 2 ] ? p + ( 60'h1 << 34 ) : p ;
      p = a [ 32 ] & b [ 3 ] ? p + ( 60'h1 << 35 ) : p ;
      p = a [ 32 ] & b [ 4 ] ? p + ( 60'h1 << 36 ) : p ;
      p = a [ 32 ] & b [ 5 ] ? p + ( 60'h1 << 37 ) : p ;
      p = a [ 32 ] & b [ 6 ] ? p + ( 60'h1 << 38 ) : p ;
      p = a [ 32 ] & b [ 7 ] ? p + ( 60'h1 << 39 ) : p ;
      p = a [ 32 ] & b [ 8 ] ? p + ( 60'h1 << 40 ) : p ;
      p = a [ 32 ] & b [ 9 ] ? p + ( 60'h1 << 41 ) : p ;
      p = a [ 32 ] & b [ 10 ] ? p + ( 60'h1 << 42 ) : p ;
      p = a [ 32 ] & b [ 11 ] ? p + ( 60'h1 << 43 ) : p ;
      p = a [ 32 ] & b [ 12 ] ? p + ( 60'h1 << 44 ) : p ;
      p = a [ 32 ] & b [ 13 ] ? p + ( 60'h1 << 45 ) : p ;
      p = a [ 32 ] & b [ 14 ] ? p + ( 60'h1 << 46 ) : p ;
      p = a [ 32 ] & b [ 15 ] ? p + ( 60'h1 << 47 ) : p ;
      p = a [ 32 ] & b [ 16 ] ? p + ( 60'h1 << 48 ) : p ;
      p = a [ 32 ] & b [ 17 ] ? p + ( 60'h1 << 49 ) : p ;
      p = a [ 32 ] & b [ 18 ] ? p + ( 60'h1 << 50 ) : p ;
      p = a [ 32 ] & b [ 19 ] ? p + ( 60'h1 << 51 ) : p ;
      p = a [ 32 ] & b [ 20 ] ? p + ( 60'h1 << 52 ) : p ;
      p = a [ 32 ] & b [ 21 ] ? p + ( 60'h1 << 53 ) : p ;
      p = a [ 32 ] & b [ 22 ] ? p + ( 60'h1 << 54 ) : p ;
      p = a [ 32 ] & b [ 23 ] ? p + ( 60'h1 << 55 ) : p ;
      p = a [ 32 ] & b [ 24 ] ? p + ( 60'h1 << 56 ) : p ;
      p = a [ 32 ] & b [ 25 ] ? p + ( 60'h1 << 57 ) : p ;
      p = a [ 32 ] & b [ 26 ] ? p + ( 60'h1 << 58 ) : p ;
      p = a [ 32 ] & b [ 27 ] ? p + ( 60'h1 << 59 ) : p ;

// Bit by Bit Multiply & Divide + Modulus
// Copyright © 2022 by Gregory Scott Callen
// All Rights Reserved.

      p = a [ 33 ] & b [ 0 ] ? p + ( 60'h1 << 33 ) : p ;
      p = a [ 33 ] & b [ 1 ] ? p + ( 60'h1 << 34 ) : p ;
      p = a [ 33 ] & b [ 2 ] ? p + ( 60'h1 << 35 ) : p ;
      p = a [ 33 ] & b [ 3 ] ? p + ( 60'h1 << 36 ) : p ;
      p = a [ 33 ] & b [ 4 ] ? p + ( 60'h1 << 37 ) : p ;
      p = a [ 33 ] & b [ 5 ] ? p + ( 60'h1 << 38 ) : p ;
      p = a [ 33 ] & b [ 6 ] ? p + ( 60'h1 << 39 ) : p ;
      p = a [ 33 ] & b [ 7 ] ? p + ( 60'h1 << 40 ) : p ;
      p = a [ 33 ] & b [ 8 ] ? p + ( 60'h1 << 41 ) : p ;
      p = a [ 33 ] & b [ 9 ] ? p + ( 60'h1 << 42 ) : p ;
      p = a [ 33 ] & b [ 10 ] ? p + ( 60'h1 << 43 ) : p ;
      p = a [ 33 ] & b [ 11 ] ? p + ( 60'h1 << 44 ) : p ;
      p = a [ 33 ] & b [ 12 ] ? p + ( 60'h1 << 45 ) : p ;
      p = a [ 33 ] & b [ 13 ] ? p + ( 60'h1 << 46 ) : p ;
      p = a [ 33 ] & b [ 14 ] ? p + ( 60'h1 << 47 ) : p ;
      p = a [ 33 ] & b [ 15 ] ? p + ( 60'h1 << 48 ) : p ;
      p = a [ 33 ] & b [ 16 ] ? p + ( 60'h1 << 49 ) : p ;
      p = a [ 33 ] & b [ 17 ] ? p + ( 60'h1 << 50 ) : p ;
      p = a [ 33 ] & b [ 18 ] ? p + ( 60'h1 << 51 ) : p ;
      p = a [ 33 ] & b [ 19 ] ? p + ( 60'h1 << 52 ) : p ;
      p = a [ 33 ] & b [ 20 ] ? p + ( 60'h1 << 53 ) : p ;
      p = a [ 33 ] & b [ 21 ] ? p + ( 60'h1 << 54 ) : p ;
      p = a [ 33 ] & b [ 22 ] ? p + ( 60'h1 << 55 ) : p ;
      p = a [ 33 ] & b [ 23 ] ? p + ( 60'h1 << 56 ) : p ;
      p = a [ 33 ] & b [ 24 ] ? p + ( 60'h1 << 57 ) : p ;
      p = a [ 33 ] & b [ 25 ] ? p + ( 60'h1 << 58 ) : p ;
      p = a [ 33 ] & b [ 26 ] ? p + ( 60'h1 << 59 ) : p ;

// Bit by Bit Multiply & Divide + Modulus
// Copyright © 2022 by Gregory Scott Callen
// All Rights Reserved.

      p = a [ 34 ] & b [ 0 ] ? p + ( 60'h1 << 34 ) : p ;
      p = a [ 34 ] & b [ 1 ] ? p + ( 60'h1 << 35 ) : p ;
      p = a [ 34 ] & b [ 2 ] ? p + ( 60'h1 << 36 ) : p ;
      p = a [ 34 ] & b [ 3 ] ? p + ( 60'h1 << 37 ) : p ;
      p = a [ 34 ] & b [ 4 ] ? p + ( 60'h1 << 38 ) : p ;
      p = a [ 34 ] & b [ 5 ] ? p + ( 60'h1 << 39 ) : p ;
      p = a [ 34 ] & b [ 6 ] ? p + ( 60'h1 << 40 ) : p ;
      p = a [ 34 ] & b [ 7 ] ? p + ( 60'h1 << 41 ) : p ;
      p = a [ 34 ] & b [ 8 ] ? p + ( 60'h1 << 42 ) : p ;
      p = a [ 34 ] & b [ 9 ] ? p + ( 60'h1 << 43 ) : p ;
      p = a [ 34 ] & b [ 10 ] ? p + ( 60'h1 << 44 ) : p ;
      p = a [ 34 ] & b [ 11 ] ? p + ( 60'h1 << 45 ) : p ;
      p = a [ 34 ] & b [ 12 ] ? p + ( 60'h1 << 46 ) : p ;
      p = a [ 34 ] & b [ 13 ] ? p + ( 60'h1 << 47 ) : p ;
      p = a [ 34 ] & b [ 14 ] ? p + ( 60'h1 << 48 ) : p ;
      p = a [ 34 ] & b [ 15 ] ? p + ( 60'h1 << 49 ) : p ;
      p = a [ 34 ] & b [ 16 ] ? p + ( 60'h1 << 50 ) : p ;
      p = a [ 34 ] & b [ 17 ] ? p + ( 60'h1 << 51 ) : p ;
      p = a [ 34 ] & b [ 18 ] ? p + ( 60'h1 << 52 ) : p ;
      p = a [ 34 ] & b [ 19 ] ? p + ( 60'h1 << 53 ) : p ;
      p = a [ 34 ] & b [ 20 ] ? p + ( 60'h1 << 54 ) : p ;
      p = a [ 34 ] & b [ 21 ] ? p + ( 60'h1 << 55 ) : p ;
      p = a [ 34 ] & b [ 22 ] ? p + ( 60'h1 << 56 ) : p ;
      p = a [ 34 ] & b [ 23 ] ? p + ( 60'h1 << 57 ) : p ;
      p = a [ 34 ] & b [ 24 ] ? p + ( 60'h1 << 58 ) : p ;
      p = a [ 34 ] & b [ 25 ] ? p + ( 60'h1 << 59 ) : p ;

// Bit by Bit Multiply & Divide + Modulus
// Copyright © 2022 by Gregory Scott Callen
// All Rights Reserved.

      p = a [ 35 ] & b [ 0 ] ? p + ( 60'h1 << 35 ) : p ;
      p = a [ 35 ] & b [ 1 ] ? p + ( 60'h1 << 36 ) : p ;
      p = a [ 35 ] & b [ 2 ] ? p + ( 60'h1 << 37 ) : p ;
      p = a [ 35 ] & b [ 3 ] ? p + ( 60'h1 << 38 ) : p ;
      p = a [ 35 ] & b [ 4 ] ? p + ( 60'h1 << 39 ) : p ;
      p = a [ 35 ] & b [ 5 ] ? p + ( 60'h1 << 40 ) : p ;
      p = a [ 35 ] & b [ 6 ] ? p + ( 60'h1 << 41 ) : p ;
      p = a [ 35 ] & b [ 7 ] ? p + ( 60'h1 << 42 ) : p ;
      p = a [ 35 ] & b [ 8 ] ? p + ( 60'h1 << 43 ) : p ;
      p = a [ 35 ] & b [ 9 ] ? p + ( 60'h1 << 44 ) : p ;
      p = a [ 35 ] & b [ 10 ] ? p + ( 60'h1 << 45 ) : p ;
      p = a [ 35 ] & b [ 11 ] ? p + ( 60'h1 << 46 ) : p ;
      p = a [ 35 ] & b [ 12 ] ? p + ( 60'h1 << 47 ) : p ;
      p = a [ 35 ] & b [ 13 ] ? p + ( 60'h1 << 48 ) : p ;
      p = a [ 35 ] & b [ 14 ] ? p + ( 60'h1 << 49 ) : p ;
      p = a [ 35 ] & b [ 15 ] ? p + ( 60'h1 << 50 ) : p ;
      p = a [ 35 ] & b [ 16 ] ? p + ( 60'h1 << 51 ) : p ;
      p = a [ 35 ] & b [ 17 ] ? p + ( 60'h1 << 52 ) : p ;
      p = a [ 35 ] & b [ 18 ] ? p + ( 60'h1 << 53 ) : p ;
      p = a [ 35 ] & b [ 19 ] ? p + ( 60'h1 << 54 ) : p ;
      p = a [ 35 ] & b [ 20 ] ? p + ( 60'h1 << 55 ) : p ;
      p = a [ 35 ] & b [ 21 ] ? p + ( 60'h1 << 56 ) : p ;
      p = a [ 35 ] & b [ 22 ] ? p + ( 60'h1 << 57 ) : p ;
      p = a [ 35 ] & b [ 23 ] ? p + ( 60'h1 << 58 ) : p ;
      p = a [ 35 ] & b [ 24 ] ? p + ( 60'h1 << 59 ) : p ;

// Bit by Bit Multiply & Divide + Modulus
// Copyright © 2022 by Gregory Scott Callen
// All Rights Reserved.

      p = a [ 36 ] & b [ 0 ] ? p + ( 60'h1 << 36 ) : p ;
      p = a [ 36 ] & b [ 1 ] ? p + ( 60'h1 << 37 ) : p ;
      p = a [ 36 ] & b [ 2 ] ? p + ( 60'h1 << 38 ) : p ;
      p = a [ 36 ] & b [ 3 ] ? p + ( 60'h1 << 39 ) : p ;
      p = a [ 36 ] & b [ 4 ] ? p + ( 60'h1 << 40 ) : p ;
      p = a [ 36 ] & b [ 5 ] ? p + ( 60'h1 << 41 ) : p ;
      p = a [ 36 ] & b [ 6 ] ? p + ( 60'h1 << 42 ) : p ;
      p = a [ 36 ] & b [ 7 ] ? p + ( 60'h1 << 43 ) : p ;
      p = a [ 36 ] & b [ 8 ] ? p + ( 60'h1 << 44 ) : p ;
      p = a [ 36 ] & b [ 9 ] ? p + ( 60'h1 << 45 ) : p ;
      p = a [ 36 ] & b [ 10 ] ? p + ( 60'h1 << 46 ) : p ;
      p = a [ 36 ] & b [ 11 ] ? p + ( 60'h1 << 47 ) : p ;
      p = a [ 36 ] & b [ 12 ] ? p + ( 60'h1 << 48 ) : p ;
      p = a [ 36 ] & b [ 13 ] ? p + ( 60'h1 << 49 ) : p ;
      p = a [ 36 ] & b [ 14 ] ? p + ( 60'h1 << 50 ) : p ;
      p = a [ 36 ] & b [ 15 ] ? p + ( 60'h1 << 51 ) : p ;
      p = a [ 36 ] & b [ 16 ] ? p + ( 60'h1 << 52 ) : p ;
      p = a [ 36 ] & b [ 17 ] ? p + ( 60'h1 << 53 ) : p ;
      p = a [ 36 ] & b [ 18 ] ? p + ( 60'h1 << 54 ) : p ;
      p = a [ 36 ] & b [ 19 ] ? p + ( 60'h1 << 55 ) : p ;
      p = a [ 36 ] & b [ 20 ] ? p + ( 60'h1 << 56 ) : p ;
      p = a [ 36 ] & b [ 21 ] ? p + ( 60'h1 << 57 ) : p ;
      p = a [ 36 ] & b [ 22 ] ? p + ( 60'h1 << 58 ) : p ;
      p = a [ 36 ] & b [ 23 ] ? p + ( 60'h1 << 59 ) : p ;

// Bit by Bit Multiply & Divide + Modulus
// Copyright © 2022 by Gregory Scott Callen
// All Rights Reserved.

      p = a [ 37 ] & b [ 0 ] ? p + ( 60'h1 << 37 ) : p ;
      p = a [ 37 ] & b [ 1 ] ? p + ( 60'h1 << 38 ) : p ;
      p = a [ 37 ] & b [ 2 ] ? p + ( 60'h1 << 39 ) : p ;
      p = a [ 37 ] & b [ 3 ] ? p + ( 60'h1 << 40 ) : p ;
      p = a [ 37 ] & b [ 4 ] ? p + ( 60'h1 << 41 ) : p ;
      p = a [ 37 ] & b [ 5 ] ? p + ( 60'h1 << 42 ) : p ;
      p = a [ 37 ] & b [ 6 ] ? p + ( 60'h1 << 43 ) : p ;
      p = a [ 37 ] & b [ 7 ] ? p + ( 60'h1 << 44 ) : p ;
      p = a [ 37 ] & b [ 8 ] ? p + ( 60'h1 << 45 ) : p ;
      p = a [ 37 ] & b [ 9 ] ? p + ( 60'h1 << 46 ) : p ;
      p = a [ 37 ] & b [ 10 ] ? p + ( 60'h1 << 47 ) : p ;
      p = a [ 37 ] & b [ 11 ] ? p + ( 60'h1 << 48 ) : p ;
      p = a [ 37 ] & b [ 12 ] ? p + ( 60'h1 << 49 ) : p ;
      p = a [ 37 ] & b [ 13 ] ? p + ( 60'h1 << 50 ) : p ;
      p = a [ 37 ] & b [ 14 ] ? p + ( 60'h1 << 51 ) : p ;
      p = a [ 37 ] & b [ 15 ] ? p + ( 60'h1 << 52 ) : p ;
      p = a [ 37 ] & b [ 16 ] ? p + ( 60'h1 << 53 ) : p ;
      p = a [ 37 ] & b [ 17 ] ? p + ( 60'h1 << 54 ) : p ;
      p = a [ 37 ] & b [ 18 ] ? p + ( 60'h1 << 55 ) : p ;
      p = a [ 37 ] & b [ 19 ] ? p + ( 60'h1 << 56 ) : p ;
      p = a [ 37 ] & b [ 20 ] ? p + ( 60'h1 << 57 ) : p ;
      p = a [ 37 ] & b [ 21 ] ? p + ( 60'h1 << 58 ) : p ;
      p = a [ 37 ] & b [ 22 ] ? p + ( 60'h1 << 59 ) : p ;

// Bit by Bit Multiply & Divide + Modulus
// Copyright © 2022 by Gregory Scott Callen
// All Rights Reserved.

      p = a [ 38 ] & b [ 0 ] ? p + ( 60'h1 << 38 ) : p ;
      p = a [ 38 ] & b [ 1 ] ? p + ( 60'h1 << 39 ) : p ;
      p = a [ 38 ] & b [ 2 ] ? p + ( 60'h1 << 40 ) : p ;
      p = a [ 38 ] & b [ 3 ] ? p + ( 60'h1 << 41 ) : p ;
      p = a [ 38 ] & b [ 4 ] ? p + ( 60'h1 << 42 ) : p ;
      p = a [ 38 ] & b [ 5 ] ? p + ( 60'h1 << 43 ) : p ;
      p = a [ 38 ] & b [ 6 ] ? p + ( 60'h1 << 44 ) : p ;
      p = a [ 38 ] & b [ 7 ] ? p + ( 60'h1 << 45 ) : p ;
      p = a [ 38 ] & b [ 8 ] ? p + ( 60'h1 << 46 ) : p ;
      p = a [ 38 ] & b [ 9 ] ? p + ( 60'h1 << 47 ) : p ;
      p = a [ 38 ] & b [ 10 ] ? p + ( 60'h1 << 48 ) : p ;
      p = a [ 38 ] & b [ 11 ] ? p + ( 60'h1 << 49 ) : p ;
      p = a [ 38 ] & b [ 12 ] ? p + ( 60'h1 << 50 ) : p ;
      p = a [ 38 ] & b [ 13 ] ? p + ( 60'h1 << 51 ) : p ;
      p = a [ 38 ] & b [ 14 ] ? p + ( 60'h1 << 52 ) : p ;
      p = a [ 38 ] & b [ 15 ] ? p + ( 60'h1 << 53 ) : p ;
      p = a [ 38 ] & b [ 16 ] ? p + ( 60'h1 << 54 ) : p ;
      p = a [ 38 ] & b [ 17 ] ? p + ( 60'h1 << 55 ) : p ;
      p = a [ 38 ] & b [ 18 ] ? p + ( 60'h1 << 56 ) : p ;
      p = a [ 38 ] & b [ 19 ] ? p + ( 60'h1 << 57 ) : p ;
      p = a [ 38 ] & b [ 20 ] ? p + ( 60'h1 << 58 ) : p ;
      p = a [ 38 ] & b [ 21 ] ? p + ( 60'h1 << 59 ) : p ;

// Bit by Bit Multiply & Divide + Modulus
// Copyright © 2022 by Gregory Scott Callen
// All Rights Reserved.

      p = a [ 39 ] & b [ 0 ] ? p + ( 60'h1 << 39 ) : p ;
      p = a [ 39 ] & b [ 1 ] ? p + ( 60'h1 << 40 ) : p ;
      p = a [ 39 ] & b [ 2 ] ? p + ( 60'h1 << 41 ) : p ;
      p = a [ 39 ] & b [ 3 ] ? p + ( 60'h1 << 42 ) : p ;
      p = a [ 39 ] & b [ 4 ] ? p + ( 60'h1 << 43 ) : p ;
      p = a [ 39 ] & b [ 5 ] ? p + ( 60'h1 << 44 ) : p ;
      p = a [ 39 ] & b [ 6 ] ? p + ( 60'h1 << 45 ) : p ;
      p = a [ 39 ] & b [ 7 ] ? p + ( 60'h1 << 46 ) : p ;
      p = a [ 39 ] & b [ 8 ] ? p + ( 60'h1 << 47 ) : p ;
      p = a [ 39 ] & b [ 9 ] ? p + ( 60'h1 << 48 ) : p ;
      p = a [ 39 ] & b [ 10 ] ? p + ( 60'h1 << 49 ) : p ;
      p = a [ 39 ] & b [ 11 ] ? p + ( 60'h1 << 50 ) : p ;
      p = a [ 39 ] & b [ 12 ] ? p + ( 60'h1 << 51 ) : p ;
      p = a [ 39 ] & b [ 13 ] ? p + ( 60'h1 << 52 ) : p ;
      p = a [ 39 ] & b [ 14 ] ? p + ( 60'h1 << 53 ) : p ;
      p = a [ 39 ] & b [ 15 ] ? p + ( 60'h1 << 54 ) : p ;
      p = a [ 39 ] & b [ 16 ] ? p + ( 60'h1 << 55 ) : p ;
      p = a [ 39 ] & b [ 17 ] ? p + ( 60'h1 << 56 ) : p ;
      p = a [ 39 ] & b [ 18 ] ? p + ( 60'h1 << 57 ) : p ;
      p = a [ 39 ] & b [ 19 ] ? p + ( 60'h1 << 58 ) : p ;
      p = a [ 39 ] & b [ 20 ] ? p + ( 60'h1 << 59 ) : p ;

// Bit by Bit Multiply & Divide + Modulus
// Copyright © 2022 by Gregory Scott Callen
// All Rights Reserved.

      p = a [ 40 ] & b [ 0 ] ? p + ( 60'h1 << 40 ) : p ;
      p = a [ 40 ] & b [ 1 ] ? p + ( 60'h1 << 41 ) : p ;
      p = a [ 40 ] & b [ 2 ] ? p + ( 60'h1 << 42 ) : p ;
      p = a [ 40 ] & b [ 3 ] ? p + ( 60'h1 << 43 ) : p ;
      p = a [ 40 ] & b [ 4 ] ? p + ( 60'h1 << 44 ) : p ;
      p = a [ 40 ] & b [ 5 ] ? p + ( 60'h1 << 45 ) : p ;
      p = a [ 40 ] & b [ 6 ] ? p + ( 60'h1 << 46 ) : p ;
      p = a [ 40 ] & b [ 7 ] ? p + ( 60'h1 << 47 ) : p ;
      p = a [ 40 ] & b [ 8 ] ? p + ( 60'h1 << 48 ) : p ;
      p = a [ 40 ] & b [ 9 ] ? p + ( 60'h1 << 49 ) : p ;
      p = a [ 40 ] & b [ 10 ] ? p + ( 60'h1 << 50 ) : p ;
      p = a [ 40 ] & b [ 11 ] ? p + ( 60'h1 << 51 ) : p ;
      p = a [ 40 ] & b [ 12 ] ? p + ( 60'h1 << 52 ) : p ;
      p = a [ 40 ] & b [ 13 ] ? p + ( 60'h1 << 53 ) : p ;
      p = a [ 40 ] & b [ 14 ] ? p + ( 60'h1 << 54 ) : p ;
      p = a [ 40 ] & b [ 15 ] ? p + ( 60'h1 << 55 ) : p ;
      p = a [ 40 ] & b [ 16 ] ? p + ( 60'h1 << 56 ) : p ;
      p = a [ 40 ] & b [ 17 ] ? p + ( 60'h1 << 57 ) : p ;
      p = a [ 40 ] & b [ 18 ] ? p + ( 60'h1 << 58 ) : p ;
      p = a [ 40 ] & b [ 19 ] ? p + ( 60'h1 << 59 ) : p ;

// Bit by Bit Multiply & Divide + Modulus
// Copyright © 2022 by Gregory Scott Callen
// All Rights Reserved.

      p = a [ 41 ] & b [ 0 ] ? p + ( 60'h1 << 41 ) : p ;
      p = a [ 41 ] & b [ 1 ] ? p + ( 60'h1 << 42 ) : p ;
      p = a [ 41 ] & b [ 2 ] ? p + ( 60'h1 << 43 ) : p ;
      p = a [ 41 ] & b [ 3 ] ? p + ( 60'h1 << 44 ) : p ;
      p = a [ 41 ] & b [ 4 ] ? p + ( 60'h1 << 45 ) : p ;
      p = a [ 41 ] & b [ 5 ] ? p + ( 60'h1 << 46 ) : p ;
      p = a [ 41 ] & b [ 6 ] ? p + ( 60'h1 << 47 ) : p ;
      p = a [ 41 ] & b [ 7 ] ? p + ( 60'h1 << 48 ) : p ;
      p = a [ 41 ] & b [ 8 ] ? p + ( 60'h1 << 49 ) : p ;
      p = a [ 41 ] & b [ 9 ] ? p + ( 60'h1 << 50 ) : p ;
      p = a [ 41 ] & b [ 10 ] ? p + ( 60'h1 << 51 ) : p ;
      p = a [ 41 ] & b [ 11 ] ? p + ( 60'h1 << 52 ) : p ;
      p = a [ 41 ] & b [ 12 ] ? p + ( 60'h1 << 53 ) : p ;
      p = a [ 41 ] & b [ 13 ] ? p + ( 60'h1 << 54 ) : p ;
      p = a [ 41 ] & b [ 14 ] ? p + ( 60'h1 << 55 ) : p ;
      p = a [ 41 ] & b [ 15 ] ? p + ( 60'h1 << 56 ) : p ;
      p = a [ 41 ] & b [ 16 ] ? p + ( 60'h1 << 57 ) : p ;
      p = a [ 41 ] & b [ 17 ] ? p + ( 60'h1 << 58 ) : p ;
      p = a [ 41 ] & b [ 18 ] ? p + ( 60'h1 << 59 ) : p ;

// Bit by Bit Multiply & Divide + Modulus
// Copyright © 2022 by Gregory Scott Callen
// All Rights Reserved.

      p = a [ 42 ] & b [ 0 ] ? p + ( 60'h1 << 42 ) : p ;
      p = a [ 42 ] & b [ 1 ] ? p + ( 60'h1 << 43 ) : p ;
      p = a [ 42 ] & b [ 2 ] ? p + ( 60'h1 << 44 ) : p ;
      p = a [ 42 ] & b [ 3 ] ? p + ( 60'h1 << 45 ) : p ;
      p = a [ 42 ] & b [ 4 ] ? p + ( 60'h1 << 46 ) : p ;
      p = a [ 42 ] & b [ 5 ] ? p + ( 60'h1 << 47 ) : p ;
      p = a [ 42 ] & b [ 6 ] ? p + ( 60'h1 << 48 ) : p ;
      p = a [ 42 ] & b [ 7 ] ? p + ( 60'h1 << 49 ) : p ;
      p = a [ 42 ] & b [ 8 ] ? p + ( 60'h1 << 50 ) : p ;
      p = a [ 42 ] & b [ 9 ] ? p + ( 60'h1 << 51 ) : p ;
      p = a [ 42 ] & b [ 10 ] ? p + ( 60'h1 << 52 ) : p ;
      p = a [ 42 ] & b [ 11 ] ? p + ( 60'h1 << 53 ) : p ;
      p = a [ 42 ] & b [ 12 ] ? p + ( 60'h1 << 54 ) : p ;
      p = a [ 42 ] & b [ 13 ] ? p + ( 60'h1 << 55 ) : p ;
      p = a [ 42 ] & b [ 14 ] ? p + ( 60'h1 << 56 ) : p ;
      p = a [ 42 ] & b [ 15 ] ? p + ( 60'h1 << 57 ) : p ;
      p = a [ 42 ] & b [ 16 ] ? p + ( 60'h1 << 58 ) : p ;
      p = a [ 42 ] & b [ 17 ] ? p + ( 60'h1 << 59 ) : p ;

// Bit by Bit Multiply & Divide + Modulus
// Copyright © 2022 by Gregory Scott Callen
// All Rights Reserved.

      p = a [ 43 ] & b [ 0 ] ? p + ( 60'h1 << 43 ) : p ;
      p = a [ 43 ] & b [ 1 ] ? p + ( 60'h1 << 44 ) : p ;
      p = a [ 43 ] & b [ 2 ] ? p + ( 60'h1 << 45 ) : p ;
      p = a [ 43 ] & b [ 3 ] ? p + ( 60'h1 << 46 ) : p ;
      p = a [ 43 ] & b [ 4 ] ? p + ( 60'h1 << 47 ) : p ;
      p = a [ 43 ] & b [ 5 ] ? p + ( 60'h1 << 48 ) : p ;
      p = a [ 43 ] & b [ 6 ] ? p + ( 60'h1 << 49 ) : p ;
      p = a [ 43 ] & b [ 7 ] ? p + ( 60'h1 << 50 ) : p ;
      p = a [ 43 ] & b [ 8 ] ? p + ( 60'h1 << 51 ) : p ;
      p = a [ 43 ] & b [ 9 ] ? p + ( 60'h1 << 52 ) : p ;
      p = a [ 43 ] & b [ 10 ] ? p + ( 60'h1 << 53 ) : p ;
      p = a [ 43 ] & b [ 11 ] ? p + ( 60'h1 << 54 ) : p ;
      p = a [ 43 ] & b [ 12 ] ? p + ( 60'h1 << 55 ) : p ;
      p = a [ 43 ] & b [ 13 ] ? p + ( 60'h1 << 56 ) : p ;
      p = a [ 43 ] & b [ 14 ] ? p + ( 60'h1 << 57 ) : p ;
      p = a [ 43 ] & b [ 15 ] ? p + ( 60'h1 << 58 ) : p ;
      p = a [ 43 ] & b [ 16 ] ? p + ( 60'h1 << 59 ) : p ;

// Bit by Bit Multiply & Divide + Modulus
// Copyright © 2022 by Gregory Scott Callen
// All Rights Reserved.

      p = a [ 44 ] & b [ 0 ] ? p + ( 60'h1 << 44 ) : p ;
      p = a [ 44 ] & b [ 1 ] ? p + ( 60'h1 << 45 ) : p ;
      p = a [ 44 ] & b [ 2 ] ? p + ( 60'h1 << 46 ) : p ;
      p = a [ 44 ] & b [ 3 ] ? p + ( 60'h1 << 47 ) : p ;
      p = a [ 44 ] & b [ 4 ] ? p + ( 60'h1 << 48 ) : p ;
      p = a [ 44 ] & b [ 5 ] ? p + ( 60'h1 << 49 ) : p ;
      p = a [ 44 ] & b [ 6 ] ? p + ( 60'h1 << 50 ) : p ;
      p = a [ 44 ] & b [ 7 ] ? p + ( 60'h1 << 51 ) : p ;
      p = a [ 44 ] & b [ 8 ] ? p + ( 60'h1 << 52 ) : p ;
      p = a [ 44 ] & b [ 9 ] ? p + ( 60'h1 << 53 ) : p ;
      p = a [ 44 ] & b [ 10 ] ? p + ( 60'h1 << 54 ) : p ;
      p = a [ 44 ] & b [ 11 ] ? p + ( 60'h1 << 55 ) : p ;
      p = a [ 44 ] & b [ 12 ] ? p + ( 60'h1 << 56 ) : p ;
      p = a [ 44 ] & b [ 13 ] ? p + ( 60'h1 << 57 ) : p ;
      p = a [ 44 ] & b [ 14 ] ? p + ( 60'h1 << 58 ) : p ;
      p = a [ 44 ] & b [ 15 ] ? p + ( 60'h1 << 59 ) : p ;

// Bit by Bit Multiply & Divide + Modulus
// Copyright © 2022 by Gregory Scott Callen
// All Rights Reserved.

      p = a [ 45 ] & b [ 0 ] ? p + ( 60'h1 << 45 ) : p ;
      p = a [ 45 ] & b [ 1 ] ? p + ( 60'h1 << 46 ) : p ;
      p = a [ 45 ] & b [ 2 ] ? p + ( 60'h1 << 47 ) : p ;
      p = a [ 45 ] & b [ 3 ] ? p + ( 60'h1 << 48 ) : p ;
      p = a [ 45 ] & b [ 4 ] ? p + ( 60'h1 << 49 ) : p ;
      p = a [ 45 ] & b [ 5 ] ? p + ( 60'h1 << 50 ) : p ;
      p = a [ 45 ] & b [ 6 ] ? p + ( 60'h1 << 51 ) : p ;
      p = a [ 45 ] & b [ 7 ] ? p + ( 60'h1 << 52 ) : p ;
      p = a [ 45 ] & b [ 8 ] ? p + ( 60'h1 << 53 ) : p ;
      p = a [ 45 ] & b [ 9 ] ? p + ( 60'h1 << 54 ) : p ;
      p = a [ 45 ] & b [ 10 ] ? p + ( 60'h1 << 55 ) : p ;
      p = a [ 45 ] & b [ 11 ] ? p + ( 60'h1 << 56 ) : p ;
      p = a [ 45 ] & b [ 12 ] ? p + ( 60'h1 << 57 ) : p ;
      p = a [ 45 ] & b [ 13 ] ? p + ( 60'h1 << 58 ) : p ;
      p = a [ 45 ] & b [ 14 ] ? p + ( 60'h1 << 59 ) : p ;

// Bit by Bit Multiply & Divide + Modulus
// Copyright © 2022 by Gregory Scott Callen
// All Rights Reserved.

      p = a [ 46 ] & b [ 0 ] ? p + ( 60'h1 << 46 ) : p ;
      p = a [ 46 ] & b [ 1 ] ? p + ( 60'h1 << 47 ) : p ;
      p = a [ 46 ] & b [ 2 ] ? p + ( 60'h1 << 48 ) : p ;
      p = a [ 46 ] & b [ 3 ] ? p + ( 60'h1 << 49 ) : p ;
      p = a [ 46 ] & b [ 4 ] ? p + ( 60'h1 << 50 ) : p ;
      p = a [ 46 ] & b [ 5 ] ? p + ( 60'h1 << 51 ) : p ;
      p = a [ 46 ] & b [ 6 ] ? p + ( 60'h1 << 52 ) : p ;
      p = a [ 46 ] & b [ 7 ] ? p + ( 60'h1 << 53 ) : p ;
      p = a [ 46 ] & b [ 8 ] ? p + ( 60'h1 << 54 ) : p ;
      p = a [ 46 ] & b [ 9 ] ? p + ( 60'h1 << 55 ) : p ;
      p = a [ 46 ] & b [ 10 ] ? p + ( 60'h1 << 56 ) : p ;
      p = a [ 46 ] & b [ 11 ] ? p + ( 60'h1 << 57 ) : p ;
      p = a [ 46 ] & b [ 12 ] ? p + ( 60'h1 << 58 ) : p ;
      p = a [ 46 ] & b [ 13 ] ? p + ( 60'h1 << 59 ) : p ;

// Bit by Bit Multiply & Divide + Modulus
// Copyright © 2022 by Gregory Scott Callen
// All Rights Reserved.

      p = a [ 47 ] & b [ 0 ] ? p + ( 60'h1 << 47 ) : p ;
      p = a [ 47 ] & b [ 1 ] ? p + ( 60'h1 << 48 ) : p ;
      p = a [ 47 ] & b [ 2 ] ? p + ( 60'h1 << 49 ) : p ;
      p = a [ 47 ] & b [ 3 ] ? p + ( 60'h1 << 50 ) : p ;
      p = a [ 47 ] & b [ 4 ] ? p + ( 60'h1 << 51 ) : p ;
      p = a [ 47 ] & b [ 5 ] ? p + ( 60'h1 << 52 ) : p ;
      p = a [ 47 ] & b [ 6 ] ? p + ( 60'h1 << 53 ) : p ;
      p = a [ 47 ] & b [ 7 ] ? p + ( 60'h1 << 54 ) : p ;
      p = a [ 47 ] & b [ 8 ] ? p + ( 60'h1 << 55 ) : p ;
      p = a [ 47 ] & b [ 9 ] ? p + ( 60'h1 << 56 ) : p ;
      p = a [ 47 ] & b [ 10 ] ? p + ( 60'h1 << 57 ) : p ;
      p = a [ 47 ] & b [ 11 ] ? p + ( 60'h1 << 58 ) : p ;
      p = a [ 47 ] & b [ 12 ] ? p + ( 60'h1 << 59 ) : p ;

// Bit by Bit Multiply & Divide + Modulus
// Copyright © 2022 by Gregory Scott Callen
// All Rights Reserved.

      p = a [ 48 ] & b [ 0 ] ? p + ( 60'h1 << 48 ) : p ;
      p = a [ 48 ] & b [ 1 ] ? p + ( 60'h1 << 49 ) : p ;
      p = a [ 48 ] & b [ 2 ] ? p + ( 60'h1 << 50 ) : p ;
      p = a [ 48 ] & b [ 3 ] ? p + ( 60'h1 << 51 ) : p ;
      p = a [ 48 ] & b [ 4 ] ? p + ( 60'h1 << 52 ) : p ;
      p = a [ 48 ] & b [ 5 ] ? p + ( 60'h1 << 53 ) : p ;
      p = a [ 48 ] & b [ 6 ] ? p + ( 60'h1 << 54 ) : p ;
      p = a [ 48 ] & b [ 7 ] ? p + ( 60'h1 << 55 ) : p ;
      p = a [ 48 ] & b [ 8 ] ? p + ( 60'h1 << 56 ) : p ;
      p = a [ 48 ] & b [ 9 ] ? p + ( 60'h1 << 57 ) : p ;
      p = a [ 48 ] & b [ 10 ] ? p + ( 60'h1 << 58 ) : p ;
      p = a [ 48 ] & b [ 11 ] ? p + ( 60'h1 << 59 ) : p ;

// Bit by Bit Multiply & Divide + Modulus
// Copyright © 2022 by Gregory Scott Callen
// All Rights Reserved.

      p = a [ 49 ] & b [ 0 ] ? p + ( 60'h1 << 49 ) : p ;
      p = a [ 49 ] & b [ 1 ] ? p + ( 60'h1 << 50 ) : p ;
      p = a [ 49 ] & b [ 2 ] ? p + ( 60'h1 << 51 ) : p ;
      p = a [ 49 ] & b [ 3 ] ? p + ( 60'h1 << 52 ) : p ;
      p = a [ 49 ] & b [ 4 ] ? p + ( 60'h1 << 53 ) : p ;
      p = a [ 49 ] & b [ 5 ] ? p + ( 60'h1 << 54 ) : p ;
      p = a [ 49 ] & b [ 6 ] ? p + ( 60'h1 << 55 ) : p ;
      p = a [ 49 ] & b [ 7 ] ? p + ( 60'h1 << 56 ) : p ;
      p = a [ 49 ] & b [ 8 ] ? p + ( 60'h1 << 57 ) : p ;
      p = a [ 49 ] & b [ 9 ] ? p + ( 60'h1 << 58 ) : p ;
      p = a [ 49 ] & b [ 10 ] ? p + ( 60'h1 << 59 ) : p ;

// Bit by Bit Multiply & Divide + Modulus
// Copyright © 2022 by Gregory Scott Callen
// All Rights Reserved.

      p = a [ 50 ] & b [ 0 ] ? p + ( 60'h1 << 50 ) : p ;
      p = a [ 50 ] & b [ 1 ] ? p + ( 60'h1 << 51 ) : p ;
      p = a [ 50 ] & b [ 2 ] ? p + ( 60'h1 << 52 ) : p ;
      p = a [ 50 ] & b [ 3 ] ? p + ( 60'h1 << 53 ) : p ;
      p = a [ 50 ] & b [ 4 ] ? p + ( 60'h1 << 54 ) : p ;
      p = a [ 50 ] & b [ 5 ] ? p + ( 60'h1 << 55 ) : p ;
      p = a [ 50 ] & b [ 6 ] ? p + ( 60'h1 << 56 ) : p ;
      p = a [ 50 ] & b [ 7 ] ? p + ( 60'h1 << 57 ) : p ;
      p = a [ 50 ] & b [ 8 ] ? p + ( 60'h1 << 58 ) : p ;
      p = a [ 50 ] & b [ 9 ] ? p + ( 60'h1 << 59 ) : p ;

// Bit by Bit Multiply & Divide + Modulus
// Copyright © 2022 by Gregory Scott Callen
// All Rights Reserved.

      p = a [ 51 ] & b [ 0 ] ? p + ( 60'h1 << 51 ) : p ;
      p = a [ 51 ] & b [ 1 ] ? p + ( 60'h1 << 52 ) : p ;
      p = a [ 51 ] & b [ 2 ] ? p + ( 60'h1 << 53 ) : p ;
      p = a [ 51 ] & b [ 3 ] ? p + ( 60'h1 << 54 ) : p ;
      p = a [ 51 ] & b [ 4 ] ? p + ( 60'h1 << 55 ) : p ;
      p = a [ 51 ] & b [ 5 ] ? p + ( 60'h1 << 56 ) : p ;
      p = a [ 51 ] & b [ 6 ] ? p + ( 60'h1 << 57 ) : p ;
      p = a [ 51 ] & b [ 7 ] ? p + ( 60'h1 << 58 ) : p ;
      p = a [ 51 ] & b [ 8 ] ? p + ( 60'h1 << 59 ) : p ;

// Bit by Bit Multiply & Divide + Modulus
// Copyright © 2022 by Gregory Scott Callen
// All Rights Reserved.

      p = a [ 52 ] & b [ 0 ] ? p + ( 60'h1 << 52 ) : p ;
      p = a [ 52 ] & b [ 1 ] ? p + ( 60'h1 << 53 ) : p ;
      p = a [ 52 ] & b [ 2 ] ? p + ( 60'h1 << 54 ) : p ;
      p = a [ 52 ] & b [ 3 ] ? p + ( 60'h1 << 55 ) : p ;
      p = a [ 52 ] & b [ 4 ] ? p + ( 60'h1 << 56 ) : p ;
      p = a [ 52 ] & b [ 5 ] ? p + ( 60'h1 << 57 ) : p ;
      p = a [ 52 ] & b [ 6 ] ? p + ( 60'h1 << 58 ) : p ;
      p = a [ 52 ] & b [ 7 ] ? p + ( 60'h1 << 59 ) : p ;

// Bit by Bit Multiply & Divide + Modulus
// Copyright © 2022 by Gregory Scott Callen
// All Rights Reserved.

      p = a [ 53 ] & b [ 0 ] ? p + ( 60'h1 << 53 ) : p ;
      p = a [ 53 ] & b [ 1 ] ? p + ( 60'h1 << 54 ) : p ;
      p = a [ 53 ] & b [ 2 ] ? p + ( 60'h1 << 55 ) : p ;
      p = a [ 53 ] & b [ 3 ] ? p + ( 60'h1 << 56 ) : p ;
      p = a [ 53 ] & b [ 4 ] ? p + ( 60'h1 << 57 ) : p ;
      p = a [ 53 ] & b [ 5 ] ? p + ( 60'h1 << 58 ) : p ;
      p = a [ 53 ] & b [ 6 ] ? p + ( 60'h1 << 59 ) : p ;

// Bit by Bit Multiply & Divide + Modulus
// Copyright © 2022 by Gregory Scott Callen
// All Rights Reserved.

      p = a [ 54 ] & b [ 0 ] ? p + ( 60'h1 << 54 ) : p ;
      p = a [ 54 ] & b [ 1 ] ? p + ( 60'h1 << 55 ) : p ;
      p = a [ 54 ] & b [ 2 ] ? p + ( 60'h1 << 56 ) : p ;
      p = a [ 54 ] & b [ 3 ] ? p + ( 60'h1 << 57 ) : p ;
      p = a [ 54 ] & b [ 4 ] ? p + ( 60'h1 << 58 ) : p ;
      p = a [ 54 ] & b [ 5 ] ? p + ( 60'h1 << 59 ) : p ;

// Bit by Bit Multiply & Divide + Modulus
// Copyright © 2022 by Gregory Scott Callen
// All Rights Reserved.

      p = a [ 55 ] & b [ 0 ] ? p + ( 60'h1 << 55 ) : p ;
      p = a [ 55 ] & b [ 1 ] ? p + ( 60'h1 << 56 ) : p ;
      p = a [ 55 ] & b [ 2 ] ? p + ( 60'h1 << 57 ) : p ;
      p = a [ 55 ] & b [ 3 ] ? p + ( 60'h1 << 58 ) : p ;
      p = a [ 55 ] & b [ 4 ] ? p + ( 60'h1 << 59 ) : p ;

// Bit by Bit Multiply & Divide + Modulus
// Copyright © 2022 by Gregory Scott Callen
// All Rights Reserved.

      p = a [ 56 ] & b [ 0 ] ? p + ( 60'h1 << 56 ) : p ;
      p = a [ 56 ] & b [ 1 ] ? p + ( 60'h1 << 57 ) : p ;
      p = a [ 56 ] & b [ 2 ] ? p + ( 60'h1 << 58 ) : p ;
      p = a [ 56 ] & b [ 3 ] ? p + ( 60'h1 << 59 ) : p ;

// Bit by Bit Multiply & Divide + Modulus
// Copyright © 2022 by Gregory Scott Callen
// All Rights Reserved.

      p = a [ 57 ] & b [ 0 ] ? p + ( 60'h1 << 57 ) : p ;
      p = a [ 57 ] & b [ 1 ] ? p + ( 60'h1 << 58 ) : p ;
      p = a [ 57 ] & b [ 2 ] ? p + ( 60'h1 << 59 ) : p ;

// Bit by Bit Multiply & Divide + Modulus
// Copyright © 2022 by Gregory Scott Callen
// All Rights Reserved.

      p = a [ 58 ] & b [ 0 ] ? p + ( 60'h1 << 58 ) : p ;
      p = a [ 58 ] & b [ 1 ] ? p + ( 60'h1 << 59 ) : p ;

// Bit by Bit Multiply & Divide + Modulus
// Copyright © 2022 by Gregory Scott Callen
// All Rights Reserved.

      p = a [ 59 ] & b [ 0 ] ? p + ( 60'h1 << 59 ) : p ;

// Bit by Bit Multiply & Divide + Modulus
// Copyright © 2022 by Gregory Scott Callen
// All Rights Reserved.

   end

endmodule    // 90198117197 = 639517 * 141041

// Bit by Bit Multiply & Divide + Modulus
// Copyright © 2022 by Gregory Scott Callen
// All Rights Reserved.

module div (
   input wire        t,
   input wire [59:0] a,
   input wite [59:0] b,
   output reg [59:0] n,
   output reg [59:0] r
);

   initial begin
      n = ~60'h0;
      r = ~60'h0;
   end

   always @ ( posedge t ) begin

      r = a;

      if (( b << 59n ) <= r ) begin
         n = n | 60'd576460752303423488;
         r = b [ 0 ] ? r - ( 60'd1 << 59 ) : r ;
      end

// Bit by Bit Multiply & Divide + Modulus
// Copyright © 2022 by Gregory Scott Callen
// All Rights Reserved.

      if (( b << 58n ) <= r ) begin
         n = n | 60'd288230376151711744;
         r = b [ 1 ] ? r - ( 60'd1 << 59 ) : r ;
         r = b [ 0 ] ? r - ( 60'd1 << 58 ) : r ;
      end

// Bit by Bit Multiply & Divide + Modulus
// Copyright © 2022 by Gregory Scott Callen
// All Rights Reserved.

      if (( b << 57n ) <= r ) begin
         n = n | 60'd144115188075855872;
         r = b [ 2 ] ? r - ( 60'd1 << 59 ) : r ;
         r = b [ 1 ] ? r - ( 60'd1 << 58 ) : r ;
         r = b [ 0 ] ? r - ( 60'd1 << 57 ) : r ;
      end

// Bit by Bit Multiply & Divide + Modulus
// Copyright © 2022 by Gregory Scott Callen
// All Rights Reserved.

      if (( b << 56n ) <= r ) begin
         n = n | 60'd72057594037927936;
         r = b [ 3 ] ? r - ( 60'd1 << 59 ) : r ;
         r = b [ 2 ] ? r - ( 60'd1 << 58 ) : r ;
         r = b [ 1 ] ? r - ( 60'd1 << 57 ) : r ;
         r = b [ 0 ] ? r - ( 60'd1 << 56 ) : r ;
      end

// Bit by Bit Multiply & Divide + Modulus
// Copyright © 2022 by Gregory Scott Callen
// All Rights Reserved.

      if (( b << 55n ) <= r ) begin
         n = n | 60'd36028797018963968;
         r = b [ 4 ] ? r - ( 60'd1 << 59 ) : r ;
         r = b [ 3 ] ? r - ( 60'd1 << 58 ) : r ;
         r = b [ 2 ] ? r - ( 60'd1 << 57 ) : r ;
         r = b [ 1 ] ? r - ( 60'd1 << 56 ) : r ;
         r = b [ 0 ] ? r - ( 60'd1 << 55 ) : r ;
      end

// Bit by Bit Multiply & Divide + Modulus
// Copyright © 2022 by Gregory Scott Callen
// All Rights Reserved.

      if (( b << 54n ) <= r ) begin
         n = n | 60'd18014398509481984;
         r = b [ 5 ] ? r - ( 60'd1 << 59 ) : r ;
         r = b [ 4 ] ? r - ( 60'd1 << 58 ) : r ;
         r = b [ 3 ] ? r - ( 60'd1 << 57 ) : r ;
         r = b [ 2 ] ? r - ( 60'd1 << 56 ) : r ;
         r = b [ 1 ] ? r - ( 60'd1 << 55 ) : r ;
         r = b [ 0 ] ? r - ( 60'd1 << 54 ) : r ;
      end

// Bit by Bit Multiply & Divide + Modulus
// Copyright © 2022 by Gregory Scott Callen
// All Rights Reserved.

      if (( b << 53n ) <= r ) begin
         n = n | 60'd9007199254740992;
         r = b [ 6 ] ? r - ( 60'd1 << 59 ) : r ;
         r = b [ 5 ] ? r - ( 60'd1 << 58 ) : r ;
         r = b [ 4 ] ? r - ( 60'd1 << 57 ) : r ;
         r = b [ 3 ] ? r - ( 60'd1 << 56 ) : r ;
         r = b [ 2 ] ? r - ( 60'd1 << 55 ) : r ;
         r = b [ 1 ] ? r - ( 60'd1 << 54 ) : r ;
         r = b [ 0 ] ? r - ( 60'd1 << 53 ) : r ;
      end

// Bit by Bit Multiply & Divide + Modulus
// Copyright © 2022 by Gregory Scott Callen
// All Rights Reserved.

      if (( b << 52n ) <= r ) begin
         n = n | 60'd4503599627370496;
         r = b [ 7 ] ? r - ( 60'd1 << 59 ) : r ;
         r = b [ 6 ] ? r - ( 60'd1 << 58 ) : r ;
         r = b [ 5 ] ? r - ( 60'd1 << 57 ) : r ;
         r = b [ 4 ] ? r - ( 60'd1 << 56 ) : r ;
         r = b [ 3 ] ? r - ( 60'd1 << 55 ) : r ;
         r = b [ 2 ] ? r - ( 60'd1 << 54 ) : r ;
         r = b [ 1 ] ? r - ( 60'd1 << 53 ) : r ;
         r = b [ 0 ] ? r - ( 60'd1 << 52 ) : r ;
      end

// Bit by Bit Multiply & Divide + Modulus
// Copyright © 2022 by Gregory Scott Callen
// All Rights Reserved.

      if (( b << 51n ) <= r ) begin
         n = n | 60'd2251799813685248;
         r = b [ 8 ] ? r - ( 60'd1 << 59 ) : r ;
         r = b [ 7 ] ? r - ( 60'd1 << 58 ) : r ;
         r = b [ 6 ] ? r - ( 60'd1 << 57 ) : r ;
         r = b [ 5 ] ? r - ( 60'd1 << 56 ) : r ;
         r = b [ 4 ] ? r - ( 60'd1 << 55 ) : r ;
         r = b [ 3 ] ? r - ( 60'd1 << 54 ) : r ;
         r = b [ 2 ] ? r - ( 60'd1 << 53 ) : r ;
         r = b [ 1 ] ? r - ( 60'd1 << 52 ) : r ;
         r = b [ 0 ] ? r - ( 60'd1 << 51 ) : r ;
      end

// Bit by Bit Multiply & Divide + Modulus
// Copyright © 2022 by Gregory Scott Callen
// All Rights Reserved.

      if (( b << 50n ) <= r ) begin
         n = n | 60'd1125899906842624;
         r = b [ 9 ] ? r - ( 60'd1 << 59 ) : r ;
         r = b [ 8 ] ? r - ( 60'd1 << 58 ) : r ;
         r = b [ 7 ] ? r - ( 60'd1 << 57 ) : r ;
         r = b [ 6 ] ? r - ( 60'd1 << 56 ) : r ;
         r = b [ 5 ] ? r - ( 60'd1 << 55 ) : r ;
         r = b [ 4 ] ? r - ( 60'd1 << 54 ) : r ;
         r = b [ 3 ] ? r - ( 60'd1 << 53 ) : r ;
         r = b [ 2 ] ? r - ( 60'd1 << 52 ) : r ;
         r = b [ 1 ] ? r - ( 60'd1 << 51 ) : r ;
         r = b [ 0 ] ? r - ( 60'd1 << 50 ) : r ;
      end

// Bit by Bit Multiply & Divide + Modulus
// Copyright © 2022 by Gregory Scott Callen
// All Rights Reserved.

      if (( b << 49n ) <= r ) begin
         n = n | 60'd562949953421312;
         r = b [ 10 ] ? r - ( 60'd1 << 59 ) : r ;
         r = b [ 9 ] ? r - ( 60'd1 << 58 ) : r ;
         r = b [ 8 ] ? r - ( 60'd1 << 57 ) : r ;
         r = b [ 7 ] ? r - ( 60'd1 << 56 ) : r ;
         r = b [ 6 ] ? r - ( 60'd1 << 55 ) : r ;
         r = b [ 5 ] ? r - ( 60'd1 << 54 ) : r ;
         r = b [ 4 ] ? r - ( 60'd1 << 53 ) : r ;
         r = b [ 3 ] ? r - ( 60'd1 << 52 ) : r ;
         r = b [ 2 ] ? r - ( 60'd1 << 51 ) : r ;
         r = b [ 1 ] ? r - ( 60'd1 << 50 ) : r ;
         r = b [ 0 ] ? r - ( 60'd1 << 49 ) : r ;
      end

// Bit by Bit Multiply & Divide + Modulus
// Copyright © 2022 by Gregory Scott Callen
// All Rights Reserved.

      if (( b << 48n ) <= r ) begin
         n = n | 60'd281474976710656;
         r = b [ 11 ] ? r - ( 60'd1 << 59 ) : r ;
         r = b [ 10 ] ? r - ( 60'd1 << 58 ) : r ;
         r = b [ 9 ] ? r - ( 60'd1 << 57 ) : r ;
         r = b [ 8 ] ? r - ( 60'd1 << 56 ) : r ;
         r = b [ 7 ] ? r - ( 60'd1 << 55 ) : r ;
         r = b [ 6 ] ? r - ( 60'd1 << 54 ) : r ;
         r = b [ 5 ] ? r - ( 60'd1 << 53 ) : r ;
         r = b [ 4 ] ? r - ( 60'd1 << 52 ) : r ;
         r = b [ 3 ] ? r - ( 60'd1 << 51 ) : r ;
         r = b [ 2 ] ? r - ( 60'd1 << 50 ) : r ;
         r = b [ 1 ] ? r - ( 60'd1 << 49 ) : r ;
         r = b [ 0 ] ? r - ( 60'd1 << 48 ) : r ;
      end

// Bit by Bit Multiply & Divide + Modulus
// Copyright © 2022 by Gregory Scott Callen
// All Rights Reserved.

      if (( b << 47n ) <= r ) begin
         n = n | 60'd140737488355328;
         r = b [ 12 ] ? r - ( 60'd1 << 59 ) : r ;
         r = b [ 11 ] ? r - ( 60'd1 << 58 ) : r ;
         r = b [ 10 ] ? r - ( 60'd1 << 57 ) : r ;
         r = b [ 9 ] ? r - ( 60'd1 << 56 ) : r ;
         r = b [ 8 ] ? r - ( 60'd1 << 55 ) : r ;
         r = b [ 7 ] ? r - ( 60'd1 << 54 ) : r ;
         r = b [ 6 ] ? r - ( 60'd1 << 53 ) : r ;
         r = b [ 5 ] ? r - ( 60'd1 << 52 ) : r ;
         r = b [ 4 ] ? r - ( 60'd1 << 51 ) : r ;
         r = b [ 3 ] ? r - ( 60'd1 << 50 ) : r ;
         r = b [ 2 ] ? r - ( 60'd1 << 49 ) : r ;
         r = b [ 1 ] ? r - ( 60'd1 << 48 ) : r ;
         r = b [ 0 ] ? r - ( 60'd1 << 47 ) : r ;
      end

// Bit by Bit Multiply & Divide + Modulus
// Copyright © 2022 by Gregory Scott Callen
// All Rights Reserved.

      if (( b << 46n ) <= r ) begin
         n = n | 60'd70368744177664;
         r = b [ 13 ] ? r - ( 60'd1 << 59 ) : r ;
         r = b [ 12 ] ? r - ( 60'd1 << 58 ) : r ;
         r = b [ 11 ] ? r - ( 60'd1 << 57 ) : r ;
         r = b [ 10 ] ? r - ( 60'd1 << 56 ) : r ;
         r = b [ 9 ] ? r - ( 60'd1 << 55 ) : r ;
         r = b [ 8 ] ? r - ( 60'd1 << 54 ) : r ;
         r = b [ 7 ] ? r - ( 60'd1 << 53 ) : r ;
         r = b [ 6 ] ? r - ( 60'd1 << 52 ) : r ;
         r = b [ 5 ] ? r - ( 60'd1 << 51 ) : r ;
         r = b [ 4 ] ? r - ( 60'd1 << 50 ) : r ;
         r = b [ 3 ] ? r - ( 60'd1 << 49 ) : r ;
         r = b [ 2 ] ? r - ( 60'd1 << 48 ) : r ;
         r = b [ 1 ] ? r - ( 60'd1 << 47 ) : r ;
         r = b [ 0 ] ? r - ( 60'd1 << 46 ) : r ;
      end

// Bit by Bit Multiply & Divide + Modulus
// Copyright © 2022 by Gregory Scott Callen
// All Rights Reserved.

      if (( b << 45n ) <= r ) begin
         n = n | 60'd35184372088832;
         r = b [ 14 ] ? r - ( 60'd1 << 59 ) : r ;
         r = b [ 13 ] ? r - ( 60'd1 << 58 ) : r ;
         r = b [ 12 ] ? r - ( 60'd1 << 57 ) : r ;
         r = b [ 11 ] ? r - ( 60'd1 << 56 ) : r ;
         r = b [ 10 ] ? r - ( 60'd1 << 55 ) : r ;
         r = b [ 9 ] ? r - ( 60'd1 << 54 ) : r ;
         r = b [ 8 ] ? r - ( 60'd1 << 53 ) : r ;
         r = b [ 7 ] ? r - ( 60'd1 << 52 ) : r ;
         r = b [ 6 ] ? r - ( 60'd1 << 51 ) : r ;
         r = b [ 5 ] ? r - ( 60'd1 << 50 ) : r ;
         r = b [ 4 ] ? r - ( 60'd1 << 49 ) : r ;
         r = b [ 3 ] ? r - ( 60'd1 << 48 ) : r ;
         r = b [ 2 ] ? r - ( 60'd1 << 47 ) : r ;
         r = b [ 1 ] ? r - ( 60'd1 << 46 ) : r ;
         r = b [ 0 ] ? r - ( 60'd1 << 45 ) : r ;
      end

// Bit by Bit Multiply & Divide + Modulus
// Copyright © 2022 by Gregory Scott Callen
// All Rights Reserved.

      if (( b << 44n ) <= r ) begin
         n = n | 60'd17592186044416;
         r = b [ 15 ] ? r - ( 60'd1 << 59 ) : r ;
         r = b [ 14 ] ? r - ( 60'd1 << 58 ) : r ;
         r = b [ 13 ] ? r - ( 60'd1 << 57 ) : r ;
         r = b [ 12 ] ? r - ( 60'd1 << 56 ) : r ;
         r = b [ 11 ] ? r - ( 60'd1 << 55 ) : r ;
         r = b [ 10 ] ? r - ( 60'd1 << 54 ) : r ;
         r = b [ 9 ] ? r - ( 60'd1 << 53 ) : r ;
         r = b [ 8 ] ? r - ( 60'd1 << 52 ) : r ;
         r = b [ 7 ] ? r - ( 60'd1 << 51 ) : r ;
         r = b [ 6 ] ? r - ( 60'd1 << 50 ) : r ;
         r = b [ 5 ] ? r - ( 60'd1 << 49 ) : r ;
         r = b [ 4 ] ? r - ( 60'd1 << 48 ) : r ;
         r = b [ 3 ] ? r - ( 60'd1 << 47 ) : r ;
         r = b [ 2 ] ? r - ( 60'd1 << 46 ) : r ;
         r = b [ 1 ] ? r - ( 60'd1 << 45 ) : r ;
         r = b [ 0 ] ? r - ( 60'd1 << 44 ) : r ;
      end

// Bit by Bit Multiply & Divide + Modulus
// Copyright © 2022 by Gregory Scott Callen
// All Rights Reserved.

      if (( b << 43n ) <= r ) begin
         n = n | 60'd8796093022208;
         r = b [ 16 ] ? r - ( 60'd1 << 59 ) : r ;
         r = b [ 15 ] ? r - ( 60'd1 << 58 ) : r ;
         r = b [ 14 ] ? r - ( 60'd1 << 57 ) : r ;
         r = b [ 13 ] ? r - ( 60'd1 << 56 ) : r ;
         r = b [ 12 ] ? r - ( 60'd1 << 55 ) : r ;
         r = b [ 11 ] ? r - ( 60'd1 << 54 ) : r ;
         r = b [ 10 ] ? r - ( 60'd1 << 53 ) : r ;
         r = b [ 9 ] ? r - ( 60'd1 << 52 ) : r ;
         r = b [ 8 ] ? r - ( 60'd1 << 51 ) : r ;
         r = b [ 7 ] ? r - ( 60'd1 << 50 ) : r ;
         r = b [ 6 ] ? r - ( 60'd1 << 49 ) : r ;
         r = b [ 5 ] ? r - ( 60'd1 << 48 ) : r ;
         r = b [ 4 ] ? r - ( 60'd1 << 47 ) : r ;
         r = b [ 3 ] ? r - ( 60'd1 << 46 ) : r ;
         r = b [ 2 ] ? r - ( 60'd1 << 45 ) : r ;
         r = b [ 1 ] ? r - ( 60'd1 << 44 ) : r ;
         r = b [ 0 ] ? r - ( 60'd1 << 43 ) : r ;
      end

// Bit by Bit Multiply & Divide + Modulus
// Copyright © 2022 by Gregory Scott Callen
// All Rights Reserved.

      if (( b << 42n ) <= r ) begin
         n = n | 60'd4398046511104;
         r = b [ 17 ] ? r - ( 60'd1 << 59 ) : r ;
         r = b [ 16 ] ? r - ( 60'd1 << 58 ) : r ;
         r = b [ 15 ] ? r - ( 60'd1 << 57 ) : r ;
         r = b [ 14 ] ? r - ( 60'd1 << 56 ) : r ;
         r = b [ 13 ] ? r - ( 60'd1 << 55 ) : r ;
         r = b [ 12 ] ? r - ( 60'd1 << 54 ) : r ;
         r = b [ 11 ] ? r - ( 60'd1 << 53 ) : r ;
         r = b [ 10 ] ? r - ( 60'd1 << 52 ) : r ;
         r = b [ 9 ] ? r - ( 60'd1 << 51 ) : r ;
         r = b [ 8 ] ? r - ( 60'd1 << 50 ) : r ;
         r = b [ 7 ] ? r - ( 60'd1 << 49 ) : r ;
         r = b [ 6 ] ? r - ( 60'd1 << 48 ) : r ;
         r = b [ 5 ] ? r - ( 60'd1 << 47 ) : r ;
         r = b [ 4 ] ? r - ( 60'd1 << 46 ) : r ;
         r = b [ 3 ] ? r - ( 60'd1 << 45 ) : r ;
         r = b [ 2 ] ? r - ( 60'd1 << 44 ) : r ;
         r = b [ 1 ] ? r - ( 60'd1 << 43 ) : r ;
         r = b [ 0 ] ? r - ( 60'd1 << 42 ) : r ;
      end

// Bit by Bit Multiply & Divide + Modulus
// Copyright © 2022 by Gregory Scott Callen
// All Rights Reserved.

      if (( b << 41n ) <= r ) begin
         n = n | 60'd2199023255552;
         r = b [ 18 ] ? r - ( 60'd1 << 59 ) : r ;
         r = b [ 17 ] ? r - ( 60'd1 << 58 ) : r ;
         r = b [ 16 ] ? r - ( 60'd1 << 57 ) : r ;
         r = b [ 15 ] ? r - ( 60'd1 << 56 ) : r ;
         r = b [ 14 ] ? r - ( 60'd1 << 55 ) : r ;
         r = b [ 13 ] ? r - ( 60'd1 << 54 ) : r ;
         r = b [ 12 ] ? r - ( 60'd1 << 53 ) : r ;
         r = b [ 11 ] ? r - ( 60'd1 << 52 ) : r ;
         r = b [ 10 ] ? r - ( 60'd1 << 51 ) : r ;
         r = b [ 9 ] ? r - ( 60'd1 << 50 ) : r ;
         r = b [ 8 ] ? r - ( 60'd1 << 49 ) : r ;
         r = b [ 7 ] ? r - ( 60'd1 << 48 ) : r ;
         r = b [ 6 ] ? r - ( 60'd1 << 47 ) : r ;
         r = b [ 5 ] ? r - ( 60'd1 << 46 ) : r ;
         r = b [ 4 ] ? r - ( 60'd1 << 45 ) : r ;
         r = b [ 3 ] ? r - ( 60'd1 << 44 ) : r ;
         r = b [ 2 ] ? r - ( 60'd1 << 43 ) : r ;
         r = b [ 1 ] ? r - ( 60'd1 << 42 ) : r ;
         r = b [ 0 ] ? r - ( 60'd1 << 41 ) : r ;
      end

// Bit by Bit Multiply & Divide + Modulus
// Copyright © 2022 by Gregory Scott Callen
// All Rights Reserved.

      if (( b << 40n ) <= r ) begin
         n = n | 60'd1099511627776;
         r = b [ 19 ] ? r - ( 60'd1 << 59 ) : r ;
         r = b [ 18 ] ? r - ( 60'd1 << 58 ) : r ;
         r = b [ 17 ] ? r - ( 60'd1 << 57 ) : r ;
         r = b [ 16 ] ? r - ( 60'd1 << 56 ) : r ;
         r = b [ 15 ] ? r - ( 60'd1 << 55 ) : r ;
         r = b [ 14 ] ? r - ( 60'd1 << 54 ) : r ;
         r = b [ 13 ] ? r - ( 60'd1 << 53 ) : r ;
         r = b [ 12 ] ? r - ( 60'd1 << 52 ) : r ;
         r = b [ 11 ] ? r - ( 60'd1 << 51 ) : r ;
         r = b [ 10 ] ? r - ( 60'd1 << 50 ) : r ;
         r = b [ 9 ] ? r - ( 60'd1 << 49 ) : r ;
         r = b [ 8 ] ? r - ( 60'd1 << 48 ) : r ;
         r = b [ 7 ] ? r - ( 60'd1 << 47 ) : r ;
         r = b [ 6 ] ? r - ( 60'd1 << 46 ) : r ;
         r = b [ 5 ] ? r - ( 60'd1 << 45 ) : r ;
         r = b [ 4 ] ? r - ( 60'd1 << 44 ) : r ;
         r = b [ 3 ] ? r - ( 60'd1 << 43 ) : r ;
         r = b [ 2 ] ? r - ( 60'd1 << 42 ) : r ;
         r = b [ 1 ] ? r - ( 60'd1 << 41 ) : r ;
         r = b [ 0 ] ? r - ( 60'd1 << 40 ) : r ;
      end

// Bit by Bit Multiply & Divide + Modulus
// Copyright © 2022 by Gregory Scott Callen
// All Rights Reserved.

      if (( b << 39n ) <= r ) begin
         n = n | 60'd549755813888;
         r = b [ 20 ] ? r - ( 60'd1 << 59 ) : r ;
         r = b [ 19 ] ? r - ( 60'd1 << 58 ) : r ;
         r = b [ 18 ] ? r - ( 60'd1 << 57 ) : r ;
         r = b [ 17 ] ? r - ( 60'd1 << 56 ) : r ;
         r = b [ 16 ] ? r - ( 60'd1 << 55 ) : r ;
         r = b [ 15 ] ? r - ( 60'd1 << 54 ) : r ;
         r = b [ 14 ] ? r - ( 60'd1 << 53 ) : r ;
         r = b [ 13 ] ? r - ( 60'd1 << 52 ) : r ;
         r = b [ 12 ] ? r - ( 60'd1 << 51 ) : r ;
         r = b [ 11 ] ? r - ( 60'd1 << 50 ) : r ;
         r = b [ 10 ] ? r - ( 60'd1 << 49 ) : r ;
         r = b [ 9 ] ? r - ( 60'd1 << 48 ) : r ;
         r = b [ 8 ] ? r - ( 60'd1 << 47 ) : r ;
         r = b [ 7 ] ? r - ( 60'd1 << 46 ) : r ;
         r = b [ 6 ] ? r - ( 60'd1 << 45 ) : r ;
         r = b [ 5 ] ? r - ( 60'd1 << 44 ) : r ;
         r = b [ 4 ] ? r - ( 60'd1 << 43 ) : r ;
         r = b [ 3 ] ? r - ( 60'd1 << 42 ) : r ;
         r = b [ 2 ] ? r - ( 60'd1 << 41 ) : r ;
         r = b [ 1 ] ? r - ( 60'd1 << 40 ) : r ;
         r = b [ 0 ] ? r - ( 60'd1 << 39 ) : r ;
      end

// Bit by Bit Multiply & Divide + Modulus
// Copyright © 2022 by Gregory Scott Callen
// All Rights Reserved.

      if (( b << 38n ) <= r ) begin
         n = n | 60'd274877906944;
         r = b [ 21 ] ? r - ( 60'd1 << 59 ) : r ;
         r = b [ 20 ] ? r - ( 60'd1 << 58 ) : r ;
         r = b [ 19 ] ? r - ( 60'd1 << 57 ) : r ;
         r = b [ 18 ] ? r - ( 60'd1 << 56 ) : r ;
         r = b [ 17 ] ? r - ( 60'd1 << 55 ) : r ;
         r = b [ 16 ] ? r - ( 60'd1 << 54 ) : r ;
         r = b [ 15 ] ? r - ( 60'd1 << 53 ) : r ;
         r = b [ 14 ] ? r - ( 60'd1 << 52 ) : r ;
         r = b [ 13 ] ? r - ( 60'd1 << 51 ) : r ;
         r = b [ 12 ] ? r - ( 60'd1 << 50 ) : r ;
         r = b [ 11 ] ? r - ( 60'd1 << 49 ) : r ;
         r = b [ 10 ] ? r - ( 60'd1 << 48 ) : r ;
         r = b [ 9 ] ? r - ( 60'd1 << 47 ) : r ;
         r = b [ 8 ] ? r - ( 60'd1 << 46 ) : r ;
         r = b [ 7 ] ? r - ( 60'd1 << 45 ) : r ;
         r = b [ 6 ] ? r - ( 60'd1 << 44 ) : r ;
         r = b [ 5 ] ? r - ( 60'd1 << 43 ) : r ;
         r = b [ 4 ] ? r - ( 60'd1 << 42 ) : r ;
         r = b [ 3 ] ? r - ( 60'd1 << 41 ) : r ;
         r = b [ 2 ] ? r - ( 60'd1 << 40 ) : r ;
         r = b [ 1 ] ? r - ( 60'd1 << 39 ) : r ;
         r = b [ 0 ] ? r - ( 60'd1 << 38 ) : r ;
      end

// Bit by Bit Multiply & Divide + Modulus
// Copyright © 2022 by Gregory Scott Callen
// All Rights Reserved.

      if (( b << 37n ) <= r ) begin
         n = n | 60'd137438953472;
         r = b [ 22 ] ? r - ( 60'd1 << 59 ) : r ;
         r = b [ 21 ] ? r - ( 60'd1 << 58 ) : r ;
         r = b [ 20 ] ? r - ( 60'd1 << 57 ) : r ;
         r = b [ 19 ] ? r - ( 60'd1 << 56 ) : r ;
         r = b [ 18 ] ? r - ( 60'd1 << 55 ) : r ;
         r = b [ 17 ] ? r - ( 60'd1 << 54 ) : r ;
         r = b [ 16 ] ? r - ( 60'd1 << 53 ) : r ;
         r = b [ 15 ] ? r - ( 60'd1 << 52 ) : r ;
         r = b [ 14 ] ? r - ( 60'd1 << 51 ) : r ;
         r = b [ 13 ] ? r - ( 60'd1 << 50 ) : r ;
         r = b [ 12 ] ? r - ( 60'd1 << 49 ) : r ;
         r = b [ 11 ] ? r - ( 60'd1 << 48 ) : r ;
         r = b [ 10 ] ? r - ( 60'd1 << 47 ) : r ;
         r = b [ 9 ] ? r - ( 60'd1 << 46 ) : r ;
         r = b [ 8 ] ? r - ( 60'd1 << 45 ) : r ;
         r = b [ 7 ] ? r - ( 60'd1 << 44 ) : r ;
         r = b [ 6 ] ? r - ( 60'd1 << 43 ) : r ;
         r = b [ 5 ] ? r - ( 60'd1 << 42 ) : r ;
         r = b [ 4 ] ? r - ( 60'd1 << 41 ) : r ;
         r = b [ 3 ] ? r - ( 60'd1 << 40 ) : r ;
         r = b [ 2 ] ? r - ( 60'd1 << 39 ) : r ;
         r = b [ 1 ] ? r - ( 60'd1 << 38 ) : r ;
         r = b [ 0 ] ? r - ( 60'd1 << 37 ) : r ;
      end

// Bit by Bit Multiply & Divide + Modulus
// Copyright © 2022 by Gregory Scott Callen
// All Rights Reserved.

      if (( b << 36n ) <= r ) begin
         n = n | 60'd68719476736;
         r = b [ 23 ] ? r - ( 60'd1 << 59 ) : r ;
         r = b [ 22 ] ? r - ( 60'd1 << 58 ) : r ;
         r = b [ 21 ] ? r - ( 60'd1 << 57 ) : r ;
         r = b [ 20 ] ? r - ( 60'd1 << 56 ) : r ;
         r = b [ 19 ] ? r - ( 60'd1 << 55 ) : r ;
         r = b [ 18 ] ? r - ( 60'd1 << 54 ) : r ;
         r = b [ 17 ] ? r - ( 60'd1 << 53 ) : r ;
         r = b [ 16 ] ? r - ( 60'd1 << 52 ) : r ;
         r = b [ 15 ] ? r - ( 60'd1 << 51 ) : r ;
         r = b [ 14 ] ? r - ( 60'd1 << 50 ) : r ;
         r = b [ 13 ] ? r - ( 60'd1 << 49 ) : r ;
         r = b [ 12 ] ? r - ( 60'd1 << 48 ) : r ;
         r = b [ 11 ] ? r - ( 60'd1 << 47 ) : r ;
         r = b [ 10 ] ? r - ( 60'd1 << 46 ) : r ;
         r = b [ 9 ] ? r - ( 60'd1 << 45 ) : r ;
         r = b [ 8 ] ? r - ( 60'd1 << 44 ) : r ;
         r = b [ 7 ] ? r - ( 60'd1 << 43 ) : r ;
         r = b [ 6 ] ? r - ( 60'd1 << 42 ) : r ;
         r = b [ 5 ] ? r - ( 60'd1 << 41 ) : r ;
         r = b [ 4 ] ? r - ( 60'd1 << 40 ) : r ;
         r = b [ 3 ] ? r - ( 60'd1 << 39 ) : r ;
         r = b [ 2 ] ? r - ( 60'd1 << 38 ) : r ;
         r = b [ 1 ] ? r - ( 60'd1 << 37 ) : r ;
         r = b [ 0 ] ? r - ( 60'd1 << 36 ) : r ;
      end

// Bit by Bit Multiply & Divide + Modulus
// Copyright © 2022 by Gregory Scott Callen
// All Rights Reserved.

      if (( b << 35n ) <= r ) begin
         n = n | 60'd34359738368;
         r = b [ 24 ] ? r - ( 60'd1 << 59 ) : r ;
         r = b [ 23 ] ? r - ( 60'd1 << 58 ) : r ;
         r = b [ 22 ] ? r - ( 60'd1 << 57 ) : r ;
         r = b [ 21 ] ? r - ( 60'd1 << 56 ) : r ;
         r = b [ 20 ] ? r - ( 60'd1 << 55 ) : r ;
         r = b [ 19 ] ? r - ( 60'd1 << 54 ) : r ;
         r = b [ 18 ] ? r - ( 60'd1 << 53 ) : r ;
         r = b [ 17 ] ? r - ( 60'd1 << 52 ) : r ;
         r = b [ 16 ] ? r - ( 60'd1 << 51 ) : r ;
         r = b [ 15 ] ? r - ( 60'd1 << 50 ) : r ;
         r = b [ 14 ] ? r - ( 60'd1 << 49 ) : r ;
         r = b [ 13 ] ? r - ( 60'd1 << 48 ) : r ;
         r = b [ 12 ] ? r - ( 60'd1 << 47 ) : r ;
         r = b [ 11 ] ? r - ( 60'd1 << 46 ) : r ;
         r = b [ 10 ] ? r - ( 60'd1 << 45 ) : r ;
         r = b [ 9 ] ? r - ( 60'd1 << 44 ) : r ;
         r = b [ 8 ] ? r - ( 60'd1 << 43 ) : r ;
         r = b [ 7 ] ? r - ( 60'd1 << 42 ) : r ;
         r = b [ 6 ] ? r - ( 60'd1 << 41 ) : r ;
         r = b [ 5 ] ? r - ( 60'd1 << 40 ) : r ;
         r = b [ 4 ] ? r - ( 60'd1 << 39 ) : r ;
         r = b [ 3 ] ? r - ( 60'd1 << 38 ) : r ;
         r = b [ 2 ] ? r - ( 60'd1 << 37 ) : r ;
         r = b [ 1 ] ? r - ( 60'd1 << 36 ) : r ;
         r = b [ 0 ] ? r - ( 60'd1 << 35 ) : r ;
      end

// Bit by Bit Multiply & Divide + Modulus
// Copyright © 2022 by Gregory Scott Callen
// All Rights Reserved.

      if (( b << 34n ) <= r ) begin
         n = n | 60'd17179869184;
         r = b [ 25 ] ? r - ( 60'd1 << 59 ) : r ;
         r = b [ 24 ] ? r - ( 60'd1 << 58 ) : r ;
         r = b [ 23 ] ? r - ( 60'd1 << 57 ) : r ;
         r = b [ 22 ] ? r - ( 60'd1 << 56 ) : r ;
         r = b [ 21 ] ? r - ( 60'd1 << 55 ) : r ;
         r = b [ 20 ] ? r - ( 60'd1 << 54 ) : r ;
         r = b [ 19 ] ? r - ( 60'd1 << 53 ) : r ;
         r = b [ 18 ] ? r - ( 60'd1 << 52 ) : r ;
         r = b [ 17 ] ? r - ( 60'd1 << 51 ) : r ;
         r = b [ 16 ] ? r - ( 60'd1 << 50 ) : r ;
         r = b [ 15 ] ? r - ( 60'd1 << 49 ) : r ;
         r = b [ 14 ] ? r - ( 60'd1 << 48 ) : r ;
         r = b [ 13 ] ? r - ( 60'd1 << 47 ) : r ;
         r = b [ 12 ] ? r - ( 60'd1 << 46 ) : r ;
         r = b [ 11 ] ? r - ( 60'd1 << 45 ) : r ;
         r = b [ 10 ] ? r - ( 60'd1 << 44 ) : r ;
         r = b [ 9 ] ? r - ( 60'd1 << 43 ) : r ;
         r = b [ 8 ] ? r - ( 60'd1 << 42 ) : r ;
         r = b [ 7 ] ? r - ( 60'd1 << 41 ) : r ;
         r = b [ 6 ] ? r - ( 60'd1 << 40 ) : r ;
         r = b [ 5 ] ? r - ( 60'd1 << 39 ) : r ;
         r = b [ 4 ] ? r - ( 60'd1 << 38 ) : r ;
         r = b [ 3 ] ? r - ( 60'd1 << 37 ) : r ;
         r = b [ 2 ] ? r - ( 60'd1 << 36 ) : r ;
         r = b [ 1 ] ? r - ( 60'd1 << 35 ) : r ;
         r = b [ 0 ] ? r - ( 60'd1 << 34 ) : r ;
      end

// Bit by Bit Multiply & Divide + Modulus
// Copyright © 2022 by Gregory Scott Callen
// All Rights Reserved.

      if (( b << 33n ) <= r ) begin
         n = n | 60'd8589934592;
         r = b [ 26 ] ? r - ( 60'd1 << 59 ) : r ;
         r = b [ 25 ] ? r - ( 60'd1 << 58 ) : r ;
         r = b [ 24 ] ? r - ( 60'd1 << 57 ) : r ;
         r = b [ 23 ] ? r - ( 60'd1 << 56 ) : r ;
         r = b [ 22 ] ? r - ( 60'd1 << 55 ) : r ;
         r = b [ 21 ] ? r - ( 60'd1 << 54 ) : r ;
         r = b [ 20 ] ? r - ( 60'd1 << 53 ) : r ;
         r = b [ 19 ] ? r - ( 60'd1 << 52 ) : r ;
         r = b [ 18 ] ? r - ( 60'd1 << 51 ) : r ;
         r = b [ 17 ] ? r - ( 60'd1 << 50 ) : r ;
         r = b [ 16 ] ? r - ( 60'd1 << 49 ) : r ;
         r = b [ 15 ] ? r - ( 60'd1 << 48 ) : r ;
         r = b [ 14 ] ? r - ( 60'd1 << 47 ) : r ;
         r = b [ 13 ] ? r - ( 60'd1 << 46 ) : r ;
         r = b [ 12 ] ? r - ( 60'd1 << 45 ) : r ;
         r = b [ 11 ] ? r - ( 60'd1 << 44 ) : r ;
         r = b [ 10 ] ? r - ( 60'd1 << 43 ) : r ;
         r = b [ 9 ] ? r - ( 60'd1 << 42 ) : r ;
         r = b [ 8 ] ? r - ( 60'd1 << 41 ) : r ;
         r = b [ 7 ] ? r - ( 60'd1 << 40 ) : r ;
         r = b [ 6 ] ? r - ( 60'd1 << 39 ) : r ;
         r = b [ 5 ] ? r - ( 60'd1 << 38 ) : r ;
         r = b [ 4 ] ? r - ( 60'd1 << 37 ) : r ;
         r = b [ 3 ] ? r - ( 60'd1 << 36 ) : r ;
         r = b [ 2 ] ? r - ( 60'd1 << 35 ) : r ;
         r = b [ 1 ] ? r - ( 60'd1 << 34 ) : r ;
         r = b [ 0 ] ? r - ( 60'd1 << 33 ) : r ;
      end

// Bit by Bit Multiply & Divide + Modulus
// Copyright © 2022 by Gregory Scott Callen
// All Rights Reserved.

      if (( b << 32n ) <= r ) begin
         n = n | 60'd4294967296;
         r = b [ 27 ] ? r - ( 60'd1 << 59 ) : r ;
         r = b [ 26 ] ? r - ( 60'd1 << 58 ) : r ;
         r = b [ 25 ] ? r - ( 60'd1 << 57 ) : r ;
         r = b [ 24 ] ? r - ( 60'd1 << 56 ) : r ;
         r = b [ 23 ] ? r - ( 60'd1 << 55 ) : r ;
         r = b [ 22 ] ? r - ( 60'd1 << 54 ) : r ;
         r = b [ 21 ] ? r - ( 60'd1 << 53 ) : r ;
         r = b [ 20 ] ? r - ( 60'd1 << 52 ) : r ;
         r = b [ 19 ] ? r - ( 60'd1 << 51 ) : r ;
         r = b [ 18 ] ? r - ( 60'd1 << 50 ) : r ;
         r = b [ 17 ] ? r - ( 60'd1 << 49 ) : r ;
         r = b [ 16 ] ? r - ( 60'd1 << 48 ) : r ;
         r = b [ 15 ] ? r - ( 60'd1 << 47 ) : r ;
         r = b [ 14 ] ? r - ( 60'd1 << 46 ) : r ;
         r = b [ 13 ] ? r - ( 60'd1 << 45 ) : r ;
         r = b [ 12 ] ? r - ( 60'd1 << 44 ) : r ;
         r = b [ 11 ] ? r - ( 60'd1 << 43 ) : r ;
         r = b [ 10 ] ? r - ( 60'd1 << 42 ) : r ;
         r = b [ 9 ] ? r - ( 60'd1 << 41 ) : r ;
         r = b [ 8 ] ? r - ( 60'd1 << 40 ) : r ;
         r = b [ 7 ] ? r - ( 60'd1 << 39 ) : r ;
         r = b [ 6 ] ? r - ( 60'd1 << 38 ) : r ;
         r = b [ 5 ] ? r - ( 60'd1 << 37 ) : r ;
         r = b [ 4 ] ? r - ( 60'd1 << 36 ) : r ;
         r = b [ 3 ] ? r - ( 60'd1 << 35 ) : r ;
         r = b [ 2 ] ? r - ( 60'd1 << 34 ) : r ;
         r = b [ 1 ] ? r - ( 60'd1 << 33 ) : r ;
         r = b [ 0 ] ? r - ( 60'd1 << 32 ) : r ;
      end

// Bit by Bit Multiply & Divide + Modulus
// Copyright © 2022 by Gregory Scott Callen
// All Rights Reserved.

      if (( b << 31n ) <= r ) begin
         n = n | 60'd2147483648;
         r = b [ 28 ] ? r - ( 60'd1 << 59 ) : r ;
         r = b [ 27 ] ? r - ( 60'd1 << 58 ) : r ;
         r = b [ 26 ] ? r - ( 60'd1 << 57 ) : r ;
         r = b [ 25 ] ? r - ( 60'd1 << 56 ) : r ;
         r = b [ 24 ] ? r - ( 60'd1 << 55 ) : r ;
         r = b [ 23 ] ? r - ( 60'd1 << 54 ) : r ;
         r = b [ 22 ] ? r - ( 60'd1 << 53 ) : r ;
         r = b [ 21 ] ? r - ( 60'd1 << 52 ) : r ;
         r = b [ 20 ] ? r - ( 60'd1 << 51 ) : r ;
         r = b [ 19 ] ? r - ( 60'd1 << 50 ) : r ;
         r = b [ 18 ] ? r - ( 60'd1 << 49 ) : r ;
         r = b [ 17 ] ? r - ( 60'd1 << 48 ) : r ;
         r = b [ 16 ] ? r - ( 60'd1 << 47 ) : r ;
         r = b [ 15 ] ? r - ( 60'd1 << 46 ) : r ;
         r = b [ 14 ] ? r - ( 60'd1 << 45 ) : r ;
         r = b [ 13 ] ? r - ( 60'd1 << 44 ) : r ;
         r = b [ 12 ] ? r - ( 60'd1 << 43 ) : r ;
         r = b [ 11 ] ? r - ( 60'd1 << 42 ) : r ;
         r = b [ 10 ] ? r - ( 60'd1 << 41 ) : r ;
         r = b [ 9 ] ? r - ( 60'd1 << 40 ) : r ;
         r = b [ 8 ] ? r - ( 60'd1 << 39 ) : r ;
         r = b [ 7 ] ? r - ( 60'd1 << 38 ) : r ;
         r = b [ 6 ] ? r - ( 60'd1 << 37 ) : r ;
         r = b [ 5 ] ? r - ( 60'd1 << 36 ) : r ;
         r = b [ 4 ] ? r - ( 60'd1 << 35 ) : r ;
         r = b [ 3 ] ? r - ( 60'd1 << 34 ) : r ;
         r = b [ 2 ] ? r - ( 60'd1 << 33 ) : r ;
         r = b [ 1 ] ? r - ( 60'd1 << 32 ) : r ;
         r = b [ 0 ] ? r - ( 60'd1 << 31 ) : r ;
      end

// Bit by Bit Multiply & Divide + Modulus
// Copyright © 2022 by Gregory Scott Callen
// All Rights Reserved.

      if (( b << 30n ) <= r ) begin
         n = n | 60'd1073741824;
         r = b [ 29 ] ? r - ( 60'd1 << 59 ) : r ;
         r = b [ 28 ] ? r - ( 60'd1 << 58 ) : r ;
         r = b [ 27 ] ? r - ( 60'd1 << 57 ) : r ;
         r = b [ 26 ] ? r - ( 60'd1 << 56 ) : r ;
         r = b [ 25 ] ? r - ( 60'd1 << 55 ) : r ;
         r = b [ 24 ] ? r - ( 60'd1 << 54 ) : r ;
         r = b [ 23 ] ? r - ( 60'd1 << 53 ) : r ;
         r = b [ 22 ] ? r - ( 60'd1 << 52 ) : r ;
         r = b [ 21 ] ? r - ( 60'd1 << 51 ) : r ;
         r = b [ 20 ] ? r - ( 60'd1 << 50 ) : r ;
         r = b [ 19 ] ? r - ( 60'd1 << 49 ) : r ;
         r = b [ 18 ] ? r - ( 60'd1 << 48 ) : r ;
         r = b [ 17 ] ? r - ( 60'd1 << 47 ) : r ;
         r = b [ 16 ] ? r - ( 60'd1 << 46 ) : r ;
         r = b [ 15 ] ? r - ( 60'd1 << 45 ) : r ;
         r = b [ 14 ] ? r - ( 60'd1 << 44 ) : r ;
         r = b [ 13 ] ? r - ( 60'd1 << 43 ) : r ;
         r = b [ 12 ] ? r - ( 60'd1 << 42 ) : r ;
         r = b [ 11 ] ? r - ( 60'd1 << 41 ) : r ;
         r = b [ 10 ] ? r - ( 60'd1 << 40 ) : r ;
         r = b [ 9 ] ? r - ( 60'd1 << 39 ) : r ;
         r = b [ 8 ] ? r - ( 60'd1 << 38 ) : r ;
         r = b [ 7 ] ? r - ( 60'd1 << 37 ) : r ;
         r = b [ 6 ] ? r - ( 60'd1 << 36 ) : r ;
         r = b [ 5 ] ? r - ( 60'd1 << 35 ) : r ;
         r = b [ 4 ] ? r - ( 60'd1 << 34 ) : r ;
         r = b [ 3 ] ? r - ( 60'd1 << 33 ) : r ;
         r = b [ 2 ] ? r - ( 60'd1 << 32 ) : r ;
         r = b [ 1 ] ? r - ( 60'd1 << 31 ) : r ;
         r = b [ 0 ] ? r - ( 60'd1 << 30 ) : r ;
      end

// Bit by Bit Multiply & Divide + Modulus
// Copyright © 2022 by Gregory Scott Callen
// All Rights Reserved.

      if (( b << 29n ) <= r ) begin
         n = n | 60'd536870912;
         r = b [ 30 ] ? r - ( 60'd1 << 59 ) : r ;
         r = b [ 29 ] ? r - ( 60'd1 << 58 ) : r ;
         r = b [ 28 ] ? r - ( 60'd1 << 57 ) : r ;
         r = b [ 27 ] ? r - ( 60'd1 << 56 ) : r ;
         r = b [ 26 ] ? r - ( 60'd1 << 55 ) : r ;
         r = b [ 25 ] ? r - ( 60'd1 << 54 ) : r ;
         r = b [ 24 ] ? r - ( 60'd1 << 53 ) : r ;
         r = b [ 23 ] ? r - ( 60'd1 << 52 ) : r ;
         r = b [ 22 ] ? r - ( 60'd1 << 51 ) : r ;
         r = b [ 21 ] ? r - ( 60'd1 << 50 ) : r ;
         r = b [ 20 ] ? r - ( 60'd1 << 49 ) : r ;
         r = b [ 19 ] ? r - ( 60'd1 << 48 ) : r ;
         r = b [ 18 ] ? r - ( 60'd1 << 47 ) : r ;
         r = b [ 17 ] ? r - ( 60'd1 << 46 ) : r ;
         r = b [ 16 ] ? r - ( 60'd1 << 45 ) : r ;
         r = b [ 15 ] ? r - ( 60'd1 << 44 ) : r ;
         r = b [ 14 ] ? r - ( 60'd1 << 43 ) : r ;
         r = b [ 13 ] ? r - ( 60'd1 << 42 ) : r ;
         r = b [ 12 ] ? r - ( 60'd1 << 41 ) : r ;
         r = b [ 11 ] ? r - ( 60'd1 << 40 ) : r ;
         r = b [ 10 ] ? r - ( 60'd1 << 39 ) : r ;
         r = b [ 9 ] ? r - ( 60'd1 << 38 ) : r ;
         r = b [ 8 ] ? r - ( 60'd1 << 37 ) : r ;
         r = b [ 7 ] ? r - ( 60'd1 << 36 ) : r ;
         r = b [ 6 ] ? r - ( 60'd1 << 35 ) : r ;
         r = b [ 5 ] ? r - ( 60'd1 << 34 ) : r ;
         r = b [ 4 ] ? r - ( 60'd1 << 33 ) : r ;
         r = b [ 3 ] ? r - ( 60'd1 << 32 ) : r ;
         r = b [ 2 ] ? r - ( 60'd1 << 31 ) : r ;
         r = b [ 1 ] ? r - ( 60'd1 << 30 ) : r ;
         r = b [ 0 ] ? r - ( 60'd1 << 29 ) : r ;
      end

// Bit by Bit Multiply & Divide + Modulus
// Copyright © 2022 by Gregory Scott Callen
// All Rights Reserved.

      if (( b << 28n ) <= r ) begin
         n = n | 60'd268435456;
         r = b [ 31 ] ? r - ( 60'd1 << 59 ) : r ;
         r = b [ 30 ] ? r - ( 60'd1 << 58 ) : r ;
         r = b [ 29 ] ? r - ( 60'd1 << 57 ) : r ;
         r = b [ 28 ] ? r - ( 60'd1 << 56 ) : r ;
         r = b [ 27 ] ? r - ( 60'd1 << 55 ) : r ;
         r = b [ 26 ] ? r - ( 60'd1 << 54 ) : r ;
         r = b [ 25 ] ? r - ( 60'd1 << 53 ) : r ;
         r = b [ 24 ] ? r - ( 60'd1 << 52 ) : r ;
         r = b [ 23 ] ? r - ( 60'd1 << 51 ) : r ;
         r = b [ 22 ] ? r - ( 60'd1 << 50 ) : r ;
         r = b [ 21 ] ? r - ( 60'd1 << 49 ) : r ;
         r = b [ 20 ] ? r - ( 60'd1 << 48 ) : r ;
         r = b [ 19 ] ? r - ( 60'd1 << 47 ) : r ;
         r = b [ 18 ] ? r - ( 60'd1 << 46 ) : r ;
         r = b [ 17 ] ? r - ( 60'd1 << 45 ) : r ;
         r = b [ 16 ] ? r - ( 60'd1 << 44 ) : r ;
         r = b [ 15 ] ? r - ( 60'd1 << 43 ) : r ;
         r = b [ 14 ] ? r - ( 60'd1 << 42 ) : r ;
         r = b [ 13 ] ? r - ( 60'd1 << 41 ) : r ;
         r = b [ 12 ] ? r - ( 60'd1 << 40 ) : r ;
         r = b [ 11 ] ? r - ( 60'd1 << 39 ) : r ;
         r = b [ 10 ] ? r - ( 60'd1 << 38 ) : r ;
         r = b [ 9 ] ? r - ( 60'd1 << 37 ) : r ;
         r = b [ 8 ] ? r - ( 60'd1 << 36 ) : r ;
         r = b [ 7 ] ? r - ( 60'd1 << 35 ) : r ;
         r = b [ 6 ] ? r - ( 60'd1 << 34 ) : r ;
         r = b [ 5 ] ? r - ( 60'd1 << 33 ) : r ;
         r = b [ 4 ] ? r - ( 60'd1 << 32 ) : r ;
         r = b [ 3 ] ? r - ( 60'd1 << 31 ) : r ;
         r = b [ 2 ] ? r - ( 60'd1 << 30 ) : r ;
         r = b [ 1 ] ? r - ( 60'd1 << 29 ) : r ;
         r = b [ 0 ] ? r - ( 60'd1 << 28 ) : r ;
      end

// Bit by Bit Multiply & Divide + Modulus
// Copyright © 2022 by Gregory Scott Callen
// All Rights Reserved.

      if (( b << 27n ) <= r ) begin
         n = n | 60'd134217728;
         r = b [ 32 ] ? r - ( 60'd1 << 59 ) : r ;
         r = b [ 31 ] ? r - ( 60'd1 << 58 ) : r ;
         r = b [ 30 ] ? r - ( 60'd1 << 57 ) : r ;
         r = b [ 29 ] ? r - ( 60'd1 << 56 ) : r ;
         r = b [ 28 ] ? r - ( 60'd1 << 55 ) : r ;
         r = b [ 27 ] ? r - ( 60'd1 << 54 ) : r ;
         r = b [ 26 ] ? r - ( 60'd1 << 53 ) : r ;
         r = b [ 25 ] ? r - ( 60'd1 << 52 ) : r ;
         r = b [ 24 ] ? r - ( 60'd1 << 51 ) : r ;
         r = b [ 23 ] ? r - ( 60'd1 << 50 ) : r ;
         r = b [ 22 ] ? r - ( 60'd1 << 49 ) : r ;
         r = b [ 21 ] ? r - ( 60'd1 << 48 ) : r ;
         r = b [ 20 ] ? r - ( 60'd1 << 47 ) : r ;
         r = b [ 19 ] ? r - ( 60'd1 << 46 ) : r ;
         r = b [ 18 ] ? r - ( 60'd1 << 45 ) : r ;
         r = b [ 17 ] ? r - ( 60'd1 << 44 ) : r ;
         r = b [ 16 ] ? r - ( 60'd1 << 43 ) : r ;
         r = b [ 15 ] ? r - ( 60'd1 << 42 ) : r ;
         r = b [ 14 ] ? r - ( 60'd1 << 41 ) : r ;
         r = b [ 13 ] ? r - ( 60'd1 << 40 ) : r ;
         r = b [ 12 ] ? r - ( 60'd1 << 39 ) : r ;
         r = b [ 11 ] ? r - ( 60'd1 << 38 ) : r ;
         r = b [ 10 ] ? r - ( 60'd1 << 37 ) : r ;
         r = b [ 9 ] ? r - ( 60'd1 << 36 ) : r ;
         r = b [ 8 ] ? r - ( 60'd1 << 35 ) : r ;
         r = b [ 7 ] ? r - ( 60'd1 << 34 ) : r ;
         r = b [ 6 ] ? r - ( 60'd1 << 33 ) : r ;
         r = b [ 5 ] ? r - ( 60'd1 << 32 ) : r ;
         r = b [ 4 ] ? r - ( 60'd1 << 31 ) : r ;
         r = b [ 3 ] ? r - ( 60'd1 << 30 ) : r ;
         r = b [ 2 ] ? r - ( 60'd1 << 29 ) : r ;
         r = b [ 1 ] ? r - ( 60'd1 << 28 ) : r ;
         r = b [ 0 ] ? r - ( 60'd1 << 27 ) : r ;
      end

// Bit by Bit Multiply & Divide + Modulus
// Copyright © 2022 by Gregory Scott Callen
// All Rights Reserved.

      if (( b << 26n ) <= r ) begin
         n = n | 60'd67108864;
         r = b [ 33 ] ? r - ( 60'd1 << 59 ) : r ;
         r = b [ 32 ] ? r - ( 60'd1 << 58 ) : r ;
         r = b [ 31 ] ? r - ( 60'd1 << 57 ) : r ;
         r = b [ 30 ] ? r - ( 60'd1 << 56 ) : r ;
         r = b [ 29 ] ? r - ( 60'd1 << 55 ) : r ;
         r = b [ 28 ] ? r - ( 60'd1 << 54 ) : r ;
         r = b [ 27 ] ? r - ( 60'd1 << 53 ) : r ;
         r = b [ 26 ] ? r - ( 60'd1 << 52 ) : r ;
         r = b [ 25 ] ? r - ( 60'd1 << 51 ) : r ;
         r = b [ 24 ] ? r - ( 60'd1 << 50 ) : r ;
         r = b [ 23 ] ? r - ( 60'd1 << 49 ) : r ;
         r = b [ 22 ] ? r - ( 60'd1 << 48 ) : r ;
         r = b [ 21 ] ? r - ( 60'd1 << 47 ) : r ;
         r = b [ 20 ] ? r - ( 60'd1 << 46 ) : r ;
         r = b [ 19 ] ? r - ( 60'd1 << 45 ) : r ;
         r = b [ 18 ] ? r - ( 60'd1 << 44 ) : r ;
         r = b [ 17 ] ? r - ( 60'd1 << 43 ) : r ;
         r = b [ 16 ] ? r - ( 60'd1 << 42 ) : r ;
         r = b [ 15 ] ? r - ( 60'd1 << 41 ) : r ;
         r = b [ 14 ] ? r - ( 60'd1 << 40 ) : r ;
         r = b [ 13 ] ? r - ( 60'd1 << 39 ) : r ;
         r = b [ 12 ] ? r - ( 60'd1 << 38 ) : r ;
         r = b [ 11 ] ? r - ( 60'd1 << 37 ) : r ;
         r = b [ 10 ] ? r - ( 60'd1 << 36 ) : r ;
         r = b [ 9 ] ? r - ( 60'd1 << 35 ) : r ;
         r = b [ 8 ] ? r - ( 60'd1 << 34 ) : r ;
         r = b [ 7 ] ? r - ( 60'd1 << 33 ) : r ;
         r = b [ 6 ] ? r - ( 60'd1 << 32 ) : r ;
         r = b [ 5 ] ? r - ( 60'd1 << 31 ) : r ;
         r = b [ 4 ] ? r - ( 60'd1 << 30 ) : r ;
         r = b [ 3 ] ? r - ( 60'd1 << 29 ) : r ;
         r = b [ 2 ] ? r - ( 60'd1 << 28 ) : r ;
         r = b [ 1 ] ? r - ( 60'd1 << 27 ) : r ;
         r = b [ 0 ] ? r - ( 60'd1 << 26 ) : r ;
      end

// Bit by Bit Multiply & Divide + Modulus
// Copyright © 2022 by Gregory Scott Callen
// All Rights Reserved.

      if (( b << 25n ) <= r ) begin
         n = n | 60'd33554432;
         r = b [ 34 ] ? r - ( 60'd1 << 59 ) : r ;
         r = b [ 33 ] ? r - ( 60'd1 << 58 ) : r ;
         r = b [ 32 ] ? r - ( 60'd1 << 57 ) : r ;
         r = b [ 31 ] ? r - ( 60'd1 << 56 ) : r ;
         r = b [ 30 ] ? r - ( 60'd1 << 55 ) : r ;
         r = b [ 29 ] ? r - ( 60'd1 << 54 ) : r ;
         r = b [ 28 ] ? r - ( 60'd1 << 53 ) : r ;
         r = b [ 27 ] ? r - ( 60'd1 << 52 ) : r ;
         r = b [ 26 ] ? r - ( 60'd1 << 51 ) : r ;
         r = b [ 25 ] ? r - ( 60'd1 << 50 ) : r ;
         r = b [ 24 ] ? r - ( 60'd1 << 49 ) : r ;
         r = b [ 23 ] ? r - ( 60'd1 << 48 ) : r ;
         r = b [ 22 ] ? r - ( 60'd1 << 47 ) : r ;
         r = b [ 21 ] ? r - ( 60'd1 << 46 ) : r ;
         r = b [ 20 ] ? r - ( 60'd1 << 45 ) : r ;
         r = b [ 19 ] ? r - ( 60'd1 << 44 ) : r ;
         r = b [ 18 ] ? r - ( 60'd1 << 43 ) : r ;
         r = b [ 17 ] ? r - ( 60'd1 << 42 ) : r ;
         r = b [ 16 ] ? r - ( 60'd1 << 41 ) : r ;
         r = b [ 15 ] ? r - ( 60'd1 << 40 ) : r ;
         r = b [ 14 ] ? r - ( 60'd1 << 39 ) : r ;
         r = b [ 13 ] ? r - ( 60'd1 << 38 ) : r ;
         r = b [ 12 ] ? r - ( 60'd1 << 37 ) : r ;
         r = b [ 11 ] ? r - ( 60'd1 << 36 ) : r ;
         r = b [ 10 ] ? r - ( 60'd1 << 35 ) : r ;
         r = b [ 9 ] ? r - ( 60'd1 << 34 ) : r ;
         r = b [ 8 ] ? r - ( 60'd1 << 33 ) : r ;
         r = b [ 7 ] ? r - ( 60'd1 << 32 ) : r ;
         r = b [ 6 ] ? r - ( 60'd1 << 31 ) : r ;
         r = b [ 5 ] ? r - ( 60'd1 << 30 ) : r ;
         r = b [ 4 ] ? r - ( 60'd1 << 29 ) : r ;
         r = b [ 3 ] ? r - ( 60'd1 << 28 ) : r ;
         r = b [ 2 ] ? r - ( 60'd1 << 27 ) : r ;
         r = b [ 1 ] ? r - ( 60'd1 << 26 ) : r ;
         r = b [ 0 ] ? r - ( 60'd1 << 25 ) : r ;
      end

// Bit by Bit Multiply & Divide + Modulus
// Copyright © 2022 by Gregory Scott Callen
// All Rights Reserved.

      if (( b << 24n ) <= r ) begin
         n = n | 60'd16777216;
         r = b [ 35 ] ? r - ( 60'd1 << 59 ) : r ;
         r = b [ 34 ] ? r - ( 60'd1 << 58 ) : r ;
         r = b [ 33 ] ? r - ( 60'd1 << 57 ) : r ;
         r = b [ 32 ] ? r - ( 60'd1 << 56 ) : r ;
         r = b [ 31 ] ? r - ( 60'd1 << 55 ) : r ;
         r = b [ 30 ] ? r - ( 60'd1 << 54 ) : r ;
         r = b [ 29 ] ? r - ( 60'd1 << 53 ) : r ;
         r = b [ 28 ] ? r - ( 60'd1 << 52 ) : r ;
         r = b [ 27 ] ? r - ( 60'd1 << 51 ) : r ;
         r = b [ 26 ] ? r - ( 60'd1 << 50 ) : r ;
         r = b [ 25 ] ? r - ( 60'd1 << 49 ) : r ;
         r = b [ 24 ] ? r - ( 60'd1 << 48 ) : r ;
         r = b [ 23 ] ? r - ( 60'd1 << 47 ) : r ;
         r = b [ 22 ] ? r - ( 60'd1 << 46 ) : r ;
         r = b [ 21 ] ? r - ( 60'd1 << 45 ) : r ;
         r = b [ 20 ] ? r - ( 60'd1 << 44 ) : r ;
         r = b [ 19 ] ? r - ( 60'd1 << 43 ) : r ;
         r = b [ 18 ] ? r - ( 60'd1 << 42 ) : r ;
         r = b [ 17 ] ? r - ( 60'd1 << 41 ) : r ;
         r = b [ 16 ] ? r - ( 60'd1 << 40 ) : r ;
         r = b [ 15 ] ? r - ( 60'd1 << 39 ) : r ;
         r = b [ 14 ] ? r - ( 60'd1 << 38 ) : r ;
         r = b [ 13 ] ? r - ( 60'd1 << 37 ) : r ;
         r = b [ 12 ] ? r - ( 60'd1 << 36 ) : r ;
         r = b [ 11 ] ? r - ( 60'd1 << 35 ) : r ;
         r = b [ 10 ] ? r - ( 60'd1 << 34 ) : r ;
         r = b [ 9 ] ? r - ( 60'd1 << 33 ) : r ;
         r = b [ 8 ] ? r - ( 60'd1 << 32 ) : r ;
         r = b [ 7 ] ? r - ( 60'd1 << 31 ) : r ;
         r = b [ 6 ] ? r - ( 60'd1 << 30 ) : r ;
         r = b [ 5 ] ? r - ( 60'd1 << 29 ) : r ;
         r = b [ 4 ] ? r - ( 60'd1 << 28 ) : r ;
         r = b [ 3 ] ? r - ( 60'd1 << 27 ) : r ;
         r = b [ 2 ] ? r - ( 60'd1 << 26 ) : r ;
         r = b [ 1 ] ? r - ( 60'd1 << 25 ) : r ;
         r = b [ 0 ] ? r - ( 60'd1 << 24 ) : r ;
      end

// Bit by Bit Multiply & Divide + Modulus
// Copyright © 2022 by Gregory Scott Callen
// All Rights Reserved.

      if (( b << 23n ) <= r ) begin
         n = n | 60'd8388608;
         r = b [ 36 ] ? r - ( 60'd1 << 59 ) : r ;
         r = b [ 35 ] ? r - ( 60'd1 << 58 ) : r ;
         r = b [ 34 ] ? r - ( 60'd1 << 57 ) : r ;
         r = b [ 33 ] ? r - ( 60'd1 << 56 ) : r ;
         r = b [ 32 ] ? r - ( 60'd1 << 55 ) : r ;
         r = b [ 31 ] ? r - ( 60'd1 << 54 ) : r ;
         r = b [ 30 ] ? r - ( 60'd1 << 53 ) : r ;
         r = b [ 29 ] ? r - ( 60'd1 << 52 ) : r ;
         r = b [ 28 ] ? r - ( 60'd1 << 51 ) : r ;
         r = b [ 27 ] ? r - ( 60'd1 << 50 ) : r ;
         r = b [ 26 ] ? r - ( 60'd1 << 49 ) : r ;
         r = b [ 25 ] ? r - ( 60'd1 << 48 ) : r ;
         r = b [ 24 ] ? r - ( 60'd1 << 47 ) : r ;
         r = b [ 23 ] ? r - ( 60'd1 << 46 ) : r ;
         r = b [ 22 ] ? r - ( 60'd1 << 45 ) : r ;
         r = b [ 21 ] ? r - ( 60'd1 << 44 ) : r ;
         r = b [ 20 ] ? r - ( 60'd1 << 43 ) : r ;
         r = b [ 19 ] ? r - ( 60'd1 << 42 ) : r ;
         r = b [ 18 ] ? r - ( 60'd1 << 41 ) : r ;
         r = b [ 17 ] ? r - ( 60'd1 << 40 ) : r ;
         r = b [ 16 ] ? r - ( 60'd1 << 39 ) : r ;
         r = b [ 15 ] ? r - ( 60'd1 << 38 ) : r ;
         r = b [ 14 ] ? r - ( 60'd1 << 37 ) : r ;
         r = b [ 13 ] ? r - ( 60'd1 << 36 ) : r ;
         r = b [ 12 ] ? r - ( 60'd1 << 35 ) : r ;
         r = b [ 11 ] ? r - ( 60'd1 << 34 ) : r ;
         r = b [ 10 ] ? r - ( 60'd1 << 33 ) : r ;
         r = b [ 9 ] ? r - ( 60'd1 << 32 ) : r ;
         r = b [ 8 ] ? r - ( 60'd1 << 31 ) : r ;
         r = b [ 7 ] ? r - ( 60'd1 << 30 ) : r ;
         r = b [ 6 ] ? r - ( 60'd1 << 29 ) : r ;
         r = b [ 5 ] ? r - ( 60'd1 << 28 ) : r ;
         r = b [ 4 ] ? r - ( 60'd1 << 27 ) : r ;
         r = b [ 3 ] ? r - ( 60'd1 << 26 ) : r ;
         r = b [ 2 ] ? r - ( 60'd1 << 25 ) : r ;
         r = b [ 1 ] ? r - ( 60'd1 << 24 ) : r ;
         r = b [ 0 ] ? r - ( 60'd1 << 23 ) : r ;
      end

// Bit by Bit Multiply & Divide + Modulus
// Copyright © 2022 by Gregory Scott Callen
// All Rights Reserved.

      if (( b << 22n ) <= r ) begin
         n = n | 60'd4194304;
         r = b [ 37 ] ? r - ( 60'd1 << 59 ) : r ;
         r = b [ 36 ] ? r - ( 60'd1 << 58 ) : r ;
         r = b [ 35 ] ? r - ( 60'd1 << 57 ) : r ;
         r = b [ 34 ] ? r - ( 60'd1 << 56 ) : r ;
         r = b [ 33 ] ? r - ( 60'd1 << 55 ) : r ;
         r = b [ 32 ] ? r - ( 60'd1 << 54 ) : r ;
         r = b [ 31 ] ? r - ( 60'd1 << 53 ) : r ;
         r = b [ 30 ] ? r - ( 60'd1 << 52 ) : r ;
         r = b [ 29 ] ? r - ( 60'd1 << 51 ) : r ;
         r = b [ 28 ] ? r - ( 60'd1 << 50 ) : r ;
         r = b [ 27 ] ? r - ( 60'd1 << 49 ) : r ;
         r = b [ 26 ] ? r - ( 60'd1 << 48 ) : r ;
         r = b [ 25 ] ? r - ( 60'd1 << 47 ) : r ;
         r = b [ 24 ] ? r - ( 60'd1 << 46 ) : r ;
         r = b [ 23 ] ? r - ( 60'd1 << 45 ) : r ;
         r = b [ 22 ] ? r - ( 60'd1 << 44 ) : r ;
         r = b [ 21 ] ? r - ( 60'd1 << 43 ) : r ;
         r = b [ 20 ] ? r - ( 60'd1 << 42 ) : r ;
         r = b [ 19 ] ? r - ( 60'd1 << 41 ) : r ;
         r = b [ 18 ] ? r - ( 60'd1 << 40 ) : r ;
         r = b [ 17 ] ? r - ( 60'd1 << 39 ) : r ;
         r = b [ 16 ] ? r - ( 60'd1 << 38 ) : r ;
         r = b [ 15 ] ? r - ( 60'd1 << 37 ) : r ;
         r = b [ 14 ] ? r - ( 60'd1 << 36 ) : r ;
         r = b [ 13 ] ? r - ( 60'd1 << 35 ) : r ;
         r = b [ 12 ] ? r - ( 60'd1 << 34 ) : r ;
         r = b [ 11 ] ? r - ( 60'd1 << 33 ) : r ;
         r = b [ 10 ] ? r - ( 60'd1 << 32 ) : r ;
         r = b [ 9 ] ? r - ( 60'd1 << 31 ) : r ;
         r = b [ 8 ] ? r - ( 60'd1 << 30 ) : r ;
         r = b [ 7 ] ? r - ( 60'd1 << 29 ) : r ;
         r = b [ 6 ] ? r - ( 60'd1 << 28 ) : r ;
         r = b [ 5 ] ? r - ( 60'd1 << 27 ) : r ;
         r = b [ 4 ] ? r - ( 60'd1 << 26 ) : r ;
         r = b [ 3 ] ? r - ( 60'd1 << 25 ) : r ;
         r = b [ 2 ] ? r - ( 60'd1 << 24 ) : r ;
         r = b [ 1 ] ? r - ( 60'd1 << 23 ) : r ;
         r = b [ 0 ] ? r - ( 60'd1 << 22 ) : r ;
      end

// Bit by Bit Multiply & Divide + Modulus
// Copyright © 2022 by Gregory Scott Callen
// All Rights Reserved.

      if (( b << 21n ) <= r ) begin
         n = n | 60'd2097152;
         r = b [ 38 ] ? r - ( 60'd1 << 59 ) : r ;
         r = b [ 37 ] ? r - ( 60'd1 << 58 ) : r ;
         r = b [ 36 ] ? r - ( 60'd1 << 57 ) : r ;
         r = b [ 35 ] ? r - ( 60'd1 << 56 ) : r ;
         r = b [ 34 ] ? r - ( 60'd1 << 55 ) : r ;
         r = b [ 33 ] ? r - ( 60'd1 << 54 ) : r ;
         r = b [ 32 ] ? r - ( 60'd1 << 53 ) : r ;
         r = b [ 31 ] ? r - ( 60'd1 << 52 ) : r ;
         r = b [ 30 ] ? r - ( 60'd1 << 51 ) : r ;
         r = b [ 29 ] ? r - ( 60'd1 << 50 ) : r ;
         r = b [ 28 ] ? r - ( 60'd1 << 49 ) : r ;
         r = b [ 27 ] ? r - ( 60'd1 << 48 ) : r ;
         r = b [ 26 ] ? r - ( 60'd1 << 47 ) : r ;
         r = b [ 25 ] ? r - ( 60'd1 << 46 ) : r ;
         r = b [ 24 ] ? r - ( 60'd1 << 45 ) : r ;
         r = b [ 23 ] ? r - ( 60'd1 << 44 ) : r ;
         r = b [ 22 ] ? r - ( 60'd1 << 43 ) : r ;
         r = b [ 21 ] ? r - ( 60'd1 << 42 ) : r ;
         r = b [ 20 ] ? r - ( 60'd1 << 41 ) : r ;
         r = b [ 19 ] ? r - ( 60'd1 << 40 ) : r ;
         r = b [ 18 ] ? r - ( 60'd1 << 39 ) : r ;
         r = b [ 17 ] ? r - ( 60'd1 << 38 ) : r ;
         r = b [ 16 ] ? r - ( 60'd1 << 37 ) : r ;
         r = b [ 15 ] ? r - ( 60'd1 << 36 ) : r ;
         r = b [ 14 ] ? r - ( 60'd1 << 35 ) : r ;
         r = b [ 13 ] ? r - ( 60'd1 << 34 ) : r ;
         r = b [ 12 ] ? r - ( 60'd1 << 33 ) : r ;
         r = b [ 11 ] ? r - ( 60'd1 << 32 ) : r ;
         r = b [ 10 ] ? r - ( 60'd1 << 31 ) : r ;
         r = b [ 9 ] ? r - ( 60'd1 << 30 ) : r ;
         r = b [ 8 ] ? r - ( 60'd1 << 29 ) : r ;
         r = b [ 7 ] ? r - ( 60'd1 << 28 ) : r ;
         r = b [ 6 ] ? r - ( 60'd1 << 27 ) : r ;
         r = b [ 5 ] ? r - ( 60'd1 << 26 ) : r ;
         r = b [ 4 ] ? r - ( 60'd1 << 25 ) : r ;
         r = b [ 3 ] ? r - ( 60'd1 << 24 ) : r ;
         r = b [ 2 ] ? r - ( 60'd1 << 23 ) : r ;
         r = b [ 1 ] ? r - ( 60'd1 << 22 ) : r ;
         r = b [ 0 ] ? r - ( 60'd1 << 21 ) : r ;
      end

// Bit by Bit Multiply & Divide + Modulus
// Copyright © 2022 by Gregory Scott Callen
// All Rights Reserved.

      if (( b << 20n ) <= r ) begin
         n = n | 60'd1048576;
         r = b [ 39 ] ? r - ( 60'd1 << 59 ) : r ;
         r = b [ 38 ] ? r - ( 60'd1 << 58 ) : r ;
         r = b [ 37 ] ? r - ( 60'd1 << 57 ) : r ;
         r = b [ 36 ] ? r - ( 60'd1 << 56 ) : r ;
         r = b [ 35 ] ? r - ( 60'd1 << 55 ) : r ;
         r = b [ 34 ] ? r - ( 60'd1 << 54 ) : r ;
         r = b [ 33 ] ? r - ( 60'd1 << 53 ) : r ;
         r = b [ 32 ] ? r - ( 60'd1 << 52 ) : r ;
         r = b [ 31 ] ? r - ( 60'd1 << 51 ) : r ;
         r = b [ 30 ] ? r - ( 60'd1 << 50 ) : r ;
         r = b [ 29 ] ? r - ( 60'd1 << 49 ) : r ;
         r = b [ 28 ] ? r - ( 60'd1 << 48 ) : r ;
         r = b [ 27 ] ? r - ( 60'd1 << 47 ) : r ;
         r = b [ 26 ] ? r - ( 60'd1 << 46 ) : r ;
         r = b [ 25 ] ? r - ( 60'd1 << 45 ) : r ;
         r = b [ 24 ] ? r - ( 60'd1 << 44 ) : r ;
         r = b [ 23 ] ? r - ( 60'd1 << 43 ) : r ;
         r = b [ 22 ] ? r - ( 60'd1 << 42 ) : r ;
         r = b [ 21 ] ? r - ( 60'd1 << 41 ) : r ;
         r = b [ 20 ] ? r - ( 60'd1 << 40 ) : r ;
         r = b [ 19 ] ? r - ( 60'd1 << 39 ) : r ;
         r = b [ 18 ] ? r - ( 60'd1 << 38 ) : r ;
         r = b [ 17 ] ? r - ( 60'd1 << 37 ) : r ;
         r = b [ 16 ] ? r - ( 60'd1 << 36 ) : r ;
         r = b [ 15 ] ? r - ( 60'd1 << 35 ) : r ;
         r = b [ 14 ] ? r - ( 60'd1 << 34 ) : r ;
         r = b [ 13 ] ? r - ( 60'd1 << 33 ) : r ;
         r = b [ 12 ] ? r - ( 60'd1 << 32 ) : r ;
         r = b [ 11 ] ? r - ( 60'd1 << 31 ) : r ;
         r = b [ 10 ] ? r - ( 60'd1 << 30 ) : r ;
         r = b [ 9 ] ? r - ( 60'd1 << 29 ) : r ;
         r = b [ 8 ] ? r - ( 60'd1 << 28 ) : r ;
         r = b [ 7 ] ? r - ( 60'd1 << 27 ) : r ;
         r = b [ 6 ] ? r - ( 60'd1 << 26 ) : r ;
         r = b [ 5 ] ? r - ( 60'd1 << 25 ) : r ;
         r = b [ 4 ] ? r - ( 60'd1 << 24 ) : r ;
         r = b [ 3 ] ? r - ( 60'd1 << 23 ) : r ;
         r = b [ 2 ] ? r - ( 60'd1 << 22 ) : r ;
         r = b [ 1 ] ? r - ( 60'd1 << 21 ) : r ;
         r = b [ 0 ] ? r - ( 60'd1 << 20 ) : r ;
      end

// Bit by Bit Multiply & Divide + Modulus
// Copyright © 2022 by Gregory Scott Callen
// All Rights Reserved.

      if (( b << 19n ) <= r ) begin
         n = n | 60'd524288;
         r = b [ 40 ] ? r - ( 60'd1 << 59 ) : r ;
         r = b [ 39 ] ? r - ( 60'd1 << 58 ) : r ;
         r = b [ 38 ] ? r - ( 60'd1 << 57 ) : r ;
         r = b [ 37 ] ? r - ( 60'd1 << 56 ) : r ;
         r = b [ 36 ] ? r - ( 60'd1 << 55 ) : r ;
         r = b [ 35 ] ? r - ( 60'd1 << 54 ) : r ;
         r = b [ 34 ] ? r - ( 60'd1 << 53 ) : r ;
         r = b [ 33 ] ? r - ( 60'd1 << 52 ) : r ;
         r = b [ 32 ] ? r - ( 60'd1 << 51 ) : r ;
         r = b [ 31 ] ? r - ( 60'd1 << 50 ) : r ;
         r = b [ 30 ] ? r - ( 60'd1 << 49 ) : r ;
         r = b [ 29 ] ? r - ( 60'd1 << 48 ) : r ;
         r = b [ 28 ] ? r - ( 60'd1 << 47 ) : r ;
         r = b [ 27 ] ? r - ( 60'd1 << 46 ) : r ;
         r = b [ 26 ] ? r - ( 60'd1 << 45 ) : r ;
         r = b [ 25 ] ? r - ( 60'd1 << 44 ) : r ;
         r = b [ 24 ] ? r - ( 60'd1 << 43 ) : r ;
         r = b [ 23 ] ? r - ( 60'd1 << 42 ) : r ;
         r = b [ 22 ] ? r - ( 60'd1 << 41 ) : r ;
         r = b [ 21 ] ? r - ( 60'd1 << 40 ) : r ;
         r = b [ 20 ] ? r - ( 60'd1 << 39 ) : r ;
         r = b [ 19 ] ? r - ( 60'd1 << 38 ) : r ;
         r = b [ 18 ] ? r - ( 60'd1 << 37 ) : r ;
         r = b [ 17 ] ? r - ( 60'd1 << 36 ) : r ;
         r = b [ 16 ] ? r - ( 60'd1 << 35 ) : r ;
         r = b [ 15 ] ? r - ( 60'd1 << 34 ) : r ;
         r = b [ 14 ] ? r - ( 60'd1 << 33 ) : r ;
         r = b [ 13 ] ? r - ( 60'd1 << 32 ) : r ;
         r = b [ 12 ] ? r - ( 60'd1 << 31 ) : r ;
         r = b [ 11 ] ? r - ( 60'd1 << 30 ) : r ;
         r = b [ 10 ] ? r - ( 60'd1 << 29 ) : r ;
         r = b [ 9 ] ? r - ( 60'd1 << 28 ) : r ;
         r = b [ 8 ] ? r - ( 60'd1 << 27 ) : r ;
         r = b [ 7 ] ? r - ( 60'd1 << 26 ) : r ;
         r = b [ 6 ] ? r - ( 60'd1 << 25 ) : r ;
         r = b [ 5 ] ? r - ( 60'd1 << 24 ) : r ;
         r = b [ 4 ] ? r - ( 60'd1 << 23 ) : r ;
         r = b [ 3 ] ? r - ( 60'd1 << 22 ) : r ;
         r = b [ 2 ] ? r - ( 60'd1 << 21 ) : r ;
         r = b [ 1 ] ? r - ( 60'd1 << 20 ) : r ;
         r = b [ 0 ] ? r - ( 60'd1 << 19 ) : r ;
      end

// Bit by Bit Multiply & Divide + Modulus
// Copyright © 2022 by Gregory Scott Callen
// All Rights Reserved.

      if (( b << 18n ) <= r ) begin
         n = n | 60'd262144;
         r = b [ 41 ] ? r - ( 60'd1 << 59 ) : r ;
         r = b [ 40 ] ? r - ( 60'd1 << 58 ) : r ;
         r = b [ 39 ] ? r - ( 60'd1 << 57 ) : r ;
         r = b [ 38 ] ? r - ( 60'd1 << 56 ) : r ;
         r = b [ 37 ] ? r - ( 60'd1 << 55 ) : r ;
         r = b [ 36 ] ? r - ( 60'd1 << 54 ) : r ;
         r = b [ 35 ] ? r - ( 60'd1 << 53 ) : r ;
         r = b [ 34 ] ? r - ( 60'd1 << 52 ) : r ;
         r = b [ 33 ] ? r - ( 60'd1 << 51 ) : r ;
         r = b [ 32 ] ? r - ( 60'd1 << 50 ) : r ;
         r = b [ 31 ] ? r - ( 60'd1 << 49 ) : r ;
         r = b [ 30 ] ? r - ( 60'd1 << 48 ) : r ;
         r = b [ 29 ] ? r - ( 60'd1 << 47 ) : r ;
         r = b [ 28 ] ? r - ( 60'd1 << 46 ) : r ;
         r = b [ 27 ] ? r - ( 60'd1 << 45 ) : r ;
         r = b [ 26 ] ? r - ( 60'd1 << 44 ) : r ;
         r = b [ 25 ] ? r - ( 60'd1 << 43 ) : r ;
         r = b [ 24 ] ? r - ( 60'd1 << 42 ) : r ;
         r = b [ 23 ] ? r - ( 60'd1 << 41 ) : r ;
         r = b [ 22 ] ? r - ( 60'd1 << 40 ) : r ;
         r = b [ 21 ] ? r - ( 60'd1 << 39 ) : r ;
         r = b [ 20 ] ? r - ( 60'd1 << 38 ) : r ;
         r = b [ 19 ] ? r - ( 60'd1 << 37 ) : r ;
         r = b [ 18 ] ? r - ( 60'd1 << 36 ) : r ;
         r = b [ 17 ] ? r - ( 60'd1 << 35 ) : r ;
         r = b [ 16 ] ? r - ( 60'd1 << 34 ) : r ;
         r = b [ 15 ] ? r - ( 60'd1 << 33 ) : r ;
         r = b [ 14 ] ? r - ( 60'd1 << 32 ) : r ;
         r = b [ 13 ] ? r - ( 60'd1 << 31 ) : r ;
         r = b [ 12 ] ? r - ( 60'd1 << 30 ) : r ;
         r = b [ 11 ] ? r - ( 60'd1 << 29 ) : r ;
         r = b [ 10 ] ? r - ( 60'd1 << 28 ) : r ;
         r = b [ 9 ] ? r - ( 60'd1 << 27 ) : r ;
         r = b [ 8 ] ? r - ( 60'd1 << 26 ) : r ;
         r = b [ 7 ] ? r - ( 60'd1 << 25 ) : r ;
         r = b [ 6 ] ? r - ( 60'd1 << 24 ) : r ;
         r = b [ 5 ] ? r - ( 60'd1 << 23 ) : r ;
         r = b [ 4 ] ? r - ( 60'd1 << 22 ) : r ;
         r = b [ 3 ] ? r - ( 60'd1 << 21 ) : r ;
         r = b [ 2 ] ? r - ( 60'd1 << 20 ) : r ;
         r = b [ 1 ] ? r - ( 60'd1 << 19 ) : r ;
         r = b [ 0 ] ? r - ( 60'd1 << 18 ) : r ;
      end

// Bit by Bit Multiply & Divide + Modulus
// Copyright © 2022 by Gregory Scott Callen
// All Rights Reserved.

      if (( b << 17n ) <= r ) begin
         n = n | 60'd131072;
         r = b [ 42 ] ? r - ( 60'd1 << 59 ) : r ;
         r = b [ 41 ] ? r - ( 60'd1 << 58 ) : r ;
         r = b [ 40 ] ? r - ( 60'd1 << 57 ) : r ;
         r = b [ 39 ] ? r - ( 60'd1 << 56 ) : r ;
         r = b [ 38 ] ? r - ( 60'd1 << 55 ) : r ;
         r = b [ 37 ] ? r - ( 60'd1 << 54 ) : r ;
         r = b [ 36 ] ? r - ( 60'd1 << 53 ) : r ;
         r = b [ 35 ] ? r - ( 60'd1 << 52 ) : r ;
         r = b [ 34 ] ? r - ( 60'd1 << 51 ) : r ;
         r = b [ 33 ] ? r - ( 60'd1 << 50 ) : r ;
         r = b [ 32 ] ? r - ( 60'd1 << 49 ) : r ;
         r = b [ 31 ] ? r - ( 60'd1 << 48 ) : r ;
         r = b [ 30 ] ? r - ( 60'd1 << 47 ) : r ;
         r = b [ 29 ] ? r - ( 60'd1 << 46 ) : r ;
         r = b [ 28 ] ? r - ( 60'd1 << 45 ) : r ;
         r = b [ 27 ] ? r - ( 60'd1 << 44 ) : r ;
         r = b [ 26 ] ? r - ( 60'd1 << 43 ) : r ;
         r = b [ 25 ] ? r - ( 60'd1 << 42 ) : r ;
         r = b [ 24 ] ? r - ( 60'd1 << 41 ) : r ;
         r = b [ 23 ] ? r - ( 60'd1 << 40 ) : r ;
         r = b [ 22 ] ? r - ( 60'd1 << 39 ) : r ;
         r = b [ 21 ] ? r - ( 60'd1 << 38 ) : r ;
         r = b [ 20 ] ? r - ( 60'd1 << 37 ) : r ;
         r = b [ 19 ] ? r - ( 60'd1 << 36 ) : r ;
         r = b [ 18 ] ? r - ( 60'd1 << 35 ) : r ;
         r = b [ 17 ] ? r - ( 60'd1 << 34 ) : r ;
         r = b [ 16 ] ? r - ( 60'd1 << 33 ) : r ;
         r = b [ 15 ] ? r - ( 60'd1 << 32 ) : r ;
         r = b [ 14 ] ? r - ( 60'd1 << 31 ) : r ;
         r = b [ 13 ] ? r - ( 60'd1 << 30 ) : r ;
         r = b [ 12 ] ? r - ( 60'd1 << 29 ) : r ;
         r = b [ 11 ] ? r - ( 60'd1 << 28 ) : r ;
         r = b [ 10 ] ? r - ( 60'd1 << 27 ) : r ;
         r = b [ 9 ] ? r - ( 60'd1 << 26 ) : r ;
         r = b [ 8 ] ? r - ( 60'd1 << 25 ) : r ;
         r = b [ 7 ] ? r - ( 60'd1 << 24 ) : r ;
         r = b [ 6 ] ? r - ( 60'd1 << 23 ) : r ;
         r = b [ 5 ] ? r - ( 60'd1 << 22 ) : r ;
         r = b [ 4 ] ? r - ( 60'd1 << 21 ) : r ;
         r = b [ 3 ] ? r - ( 60'd1 << 20 ) : r ;
         r = b [ 2 ] ? r - ( 60'd1 << 19 ) : r ;
         r = b [ 1 ] ? r - ( 60'd1 << 18 ) : r ;
         r = b [ 0 ] ? r - ( 60'd1 << 17 ) : r ;
      end

// Bit by Bit Multiply & Divide + Modulus
// Copyright © 2022 by Gregory Scott Callen
// All Rights Reserved.

      if (( b << 16n ) <= r ) begin
         n = n | 60'd65536;
         r = b [ 43 ] ? r - ( 60'd1 << 59 ) : r ;
         r = b [ 42 ] ? r - ( 60'd1 << 58 ) : r ;
         r = b [ 41 ] ? r - ( 60'd1 << 57 ) : r ;
         r = b [ 40 ] ? r - ( 60'd1 << 56 ) : r ;
         r = b [ 39 ] ? r - ( 60'd1 << 55 ) : r ;
         r = b [ 38 ] ? r - ( 60'd1 << 54 ) : r ;
         r = b [ 37 ] ? r - ( 60'd1 << 53 ) : r ;
         r = b [ 36 ] ? r - ( 60'd1 << 52 ) : r ;
         r = b [ 35 ] ? r - ( 60'd1 << 51 ) : r ;
         r = b [ 34 ] ? r - ( 60'd1 << 50 ) : r ;
         r = b [ 33 ] ? r - ( 60'd1 << 49 ) : r ;
         r = b [ 32 ] ? r - ( 60'd1 << 48 ) : r ;
         r = b [ 31 ] ? r - ( 60'd1 << 47 ) : r ;
         r = b [ 30 ] ? r - ( 60'd1 << 46 ) : r ;
         r = b [ 29 ] ? r - ( 60'd1 << 45 ) : r ;
         r = b [ 28 ] ? r - ( 60'd1 << 44 ) : r ;
         r = b [ 27 ] ? r - ( 60'd1 << 43 ) : r ;
         r = b [ 26 ] ? r - ( 60'd1 << 42 ) : r ;
         r = b [ 25 ] ? r - ( 60'd1 << 41 ) : r ;
         r = b [ 24 ] ? r - ( 60'd1 << 40 ) : r ;
         r = b [ 23 ] ? r - ( 60'd1 << 39 ) : r ;
         r = b [ 22 ] ? r - ( 60'd1 << 38 ) : r ;
         r = b [ 21 ] ? r - ( 60'd1 << 37 ) : r ;
         r = b [ 20 ] ? r - ( 60'd1 << 36 ) : r ;
         r = b [ 19 ] ? r - ( 60'd1 << 35 ) : r ;
         r = b [ 18 ] ? r - ( 60'd1 << 34 ) : r ;
         r = b [ 17 ] ? r - ( 60'd1 << 33 ) : r ;
         r = b [ 16 ] ? r - ( 60'd1 << 32 ) : r ;
         r = b [ 15 ] ? r - ( 60'd1 << 31 ) : r ;
         r = b [ 14 ] ? r - ( 60'd1 << 30 ) : r ;
         r = b [ 13 ] ? r - ( 60'd1 << 29 ) : r ;
         r = b [ 12 ] ? r - ( 60'd1 << 28 ) : r ;
         r = b [ 11 ] ? r - ( 60'd1 << 27 ) : r ;
         r = b [ 10 ] ? r - ( 60'd1 << 26 ) : r ;
         r = b [ 9 ] ? r - ( 60'd1 << 25 ) : r ;
         r = b [ 8 ] ? r - ( 60'd1 << 24 ) : r ;
         r = b [ 7 ] ? r - ( 60'd1 << 23 ) : r ;
         r = b [ 6 ] ? r - ( 60'd1 << 22 ) : r ;
         r = b [ 5 ] ? r - ( 60'd1 << 21 ) : r ;
         r = b [ 4 ] ? r - ( 60'd1 << 20 ) : r ;
         r = b [ 3 ] ? r - ( 60'd1 << 19 ) : r ;
         r = b [ 2 ] ? r - ( 60'd1 << 18 ) : r ;
         r = b [ 1 ] ? r - ( 60'd1 << 17 ) : r ;
         r = b [ 0 ] ? r - ( 60'd1 << 16 ) : r ;
      end

// Bit by Bit Multiply & Divide + Modulus
// Copyright © 2022 by Gregory Scott Callen
// All Rights Reserved.

      if (( b << 15n ) <= r ) begin
         n = n | 60'd32768;
         r = b [ 44 ] ? r - ( 60'd1 << 59 ) : r ;
         r = b [ 43 ] ? r - ( 60'd1 << 58 ) : r ;
         r = b [ 42 ] ? r - ( 60'd1 << 57 ) : r ;
         r = b [ 41 ] ? r - ( 60'd1 << 56 ) : r ;
         r = b [ 40 ] ? r - ( 60'd1 << 55 ) : r ;
         r = b [ 39 ] ? r - ( 60'd1 << 54 ) : r ;
         r = b [ 38 ] ? r - ( 60'd1 << 53 ) : r ;
         r = b [ 37 ] ? r - ( 60'd1 << 52 ) : r ;
         r = b [ 36 ] ? r - ( 60'd1 << 51 ) : r ;
         r = b [ 35 ] ? r - ( 60'd1 << 50 ) : r ;
         r = b [ 34 ] ? r - ( 60'd1 << 49 ) : r ;
         r = b [ 33 ] ? r - ( 60'd1 << 48 ) : r ;
         r = b [ 32 ] ? r - ( 60'd1 << 47 ) : r ;
         r = b [ 31 ] ? r - ( 60'd1 << 46 ) : r ;
         r = b [ 30 ] ? r - ( 60'd1 << 45 ) : r ;
         r = b [ 29 ] ? r - ( 60'd1 << 44 ) : r ;
         r = b [ 28 ] ? r - ( 60'd1 << 43 ) : r ;
         r = b [ 27 ] ? r - ( 60'd1 << 42 ) : r ;
         r = b [ 26 ] ? r - ( 60'd1 << 41 ) : r ;
         r = b [ 25 ] ? r - ( 60'd1 << 40 ) : r ;
         r = b [ 24 ] ? r - ( 60'd1 << 39 ) : r ;
         r = b [ 23 ] ? r - ( 60'd1 << 38 ) : r ;
         r = b [ 22 ] ? r - ( 60'd1 << 37 ) : r ;
         r = b [ 21 ] ? r - ( 60'd1 << 36 ) : r ;
         r = b [ 20 ] ? r - ( 60'd1 << 35 ) : r ;
         r = b [ 19 ] ? r - ( 60'd1 << 34 ) : r ;
         r = b [ 18 ] ? r - ( 60'd1 << 33 ) : r ;
         r = b [ 17 ] ? r - ( 60'd1 << 32 ) : r ;
         r = b [ 16 ] ? r - ( 60'd1 << 31 ) : r ;
         r = b [ 15 ] ? r - ( 60'd1 << 30 ) : r ;
         r = b [ 14 ] ? r - ( 60'd1 << 29 ) : r ;
         r = b [ 13 ] ? r - ( 60'd1 << 28 ) : r ;
         r = b [ 12 ] ? r - ( 60'd1 << 27 ) : r ;
         r = b [ 11 ] ? r - ( 60'd1 << 26 ) : r ;
         r = b [ 10 ] ? r - ( 60'd1 << 25 ) : r ;
         r = b [ 9 ] ? r - ( 60'd1 << 24 ) : r ;
         r = b [ 8 ] ? r - ( 60'd1 << 23 ) : r ;
         r = b [ 7 ] ? r - ( 60'd1 << 22 ) : r ;
         r = b [ 6 ] ? r - ( 60'd1 << 21 ) : r ;
         r = b [ 5 ] ? r - ( 60'd1 << 20 ) : r ;
         r = b [ 4 ] ? r - ( 60'd1 << 19 ) : r ;
         r = b [ 3 ] ? r - ( 60'd1 << 18 ) : r ;
         r = b [ 2 ] ? r - ( 60'd1 << 17 ) : r ;
         r = b [ 1 ] ? r - ( 60'd1 << 16 ) : r ;
         r = b [ 0 ] ? r - ( 60'd1 << 15 ) : r ;
      end

// Bit by Bit Multiply & Divide + Modulus
// Copyright © 2022 by Gregory Scott Callen
// All Rights Reserved.

      if (( b << 14n ) <= r ) begin
         n = n | 60'd16384;
         r = b [ 45 ] ? r - ( 60'd1 << 59 ) : r ;
         r = b [ 44 ] ? r - ( 60'd1 << 58 ) : r ;
         r = b [ 43 ] ? r - ( 60'd1 << 57 ) : r ;
         r = b [ 42 ] ? r - ( 60'd1 << 56 ) : r ;
         r = b [ 41 ] ? r - ( 60'd1 << 55 ) : r ;
         r = b [ 40 ] ? r - ( 60'd1 << 54 ) : r ;
         r = b [ 39 ] ? r - ( 60'd1 << 53 ) : r ;
         r = b [ 38 ] ? r - ( 60'd1 << 52 ) : r ;
         r = b [ 37 ] ? r - ( 60'd1 << 51 ) : r ;
         r = b [ 36 ] ? r - ( 60'd1 << 50 ) : r ;
         r = b [ 35 ] ? r - ( 60'd1 << 49 ) : r ;
         r = b [ 34 ] ? r - ( 60'd1 << 48 ) : r ;
         r = b [ 33 ] ? r - ( 60'd1 << 47 ) : r ;
         r = b [ 32 ] ? r - ( 60'd1 << 46 ) : r ;
         r = b [ 31 ] ? r - ( 60'd1 << 45 ) : r ;
         r = b [ 30 ] ? r - ( 60'd1 << 44 ) : r ;
         r = b [ 29 ] ? r - ( 60'd1 << 43 ) : r ;
         r = b [ 28 ] ? r - ( 60'd1 << 42 ) : r ;
         r = b [ 27 ] ? r - ( 60'd1 << 41 ) : r ;
         r = b [ 26 ] ? r - ( 60'd1 << 40 ) : r ;
         r = b [ 25 ] ? r - ( 60'd1 << 39 ) : r ;
         r = b [ 24 ] ? r - ( 60'd1 << 38 ) : r ;
         r = b [ 23 ] ? r - ( 60'd1 << 37 ) : r ;
         r = b [ 22 ] ? r - ( 60'd1 << 36 ) : r ;
         r = b [ 21 ] ? r - ( 60'd1 << 35 ) : r ;
         r = b [ 20 ] ? r - ( 60'd1 << 34 ) : r ;
         r = b [ 19 ] ? r - ( 60'd1 << 33 ) : r ;
         r = b [ 18 ] ? r - ( 60'd1 << 32 ) : r ;
         r = b [ 17 ] ? r - ( 60'd1 << 31 ) : r ;
         r = b [ 16 ] ? r - ( 60'd1 << 30 ) : r ;
         r = b [ 15 ] ? r - ( 60'd1 << 29 ) : r ;
         r = b [ 14 ] ? r - ( 60'd1 << 28 ) : r ;
         r = b [ 13 ] ? r - ( 60'd1 << 27 ) : r ;
         r = b [ 12 ] ? r - ( 60'd1 << 26 ) : r ;
         r = b [ 11 ] ? r - ( 60'd1 << 25 ) : r ;
         r = b [ 10 ] ? r - ( 60'd1 << 24 ) : r ;
         r = b [ 9 ] ? r - ( 60'd1 << 23 ) : r ;
         r = b [ 8 ] ? r - ( 60'd1 << 22 ) : r ;
         r = b [ 7 ] ? r - ( 60'd1 << 21 ) : r ;
         r = b [ 6 ] ? r - ( 60'd1 << 20 ) : r ;
         r = b [ 5 ] ? r - ( 60'd1 << 19 ) : r ;
         r = b [ 4 ] ? r - ( 60'd1 << 18 ) : r ;
         r = b [ 3 ] ? r - ( 60'd1 << 17 ) : r ;
         r = b [ 2 ] ? r - ( 60'd1 << 16 ) : r ;
         r = b [ 1 ] ? r - ( 60'd1 << 15 ) : r ;
         r = b [ 0 ] ? r - ( 60'd1 << 14 ) : r ;
      end

// Bit by Bit Multiply & Divide + Modulus
// Copyright © 2022 by Gregory Scott Callen
// All Rights Reserved.

      if (( b << 13n ) <= r ) begin
         n = n | 60'd8192;
         r = b [ 46 ] ? r - ( 60'd1 << 59 ) : r ;
         r = b [ 45 ] ? r - ( 60'd1 << 58 ) : r ;
         r = b [ 44 ] ? r - ( 60'd1 << 57 ) : r ;
         r = b [ 43 ] ? r - ( 60'd1 << 56 ) : r ;
         r = b [ 42 ] ? r - ( 60'd1 << 55 ) : r ;
         r = b [ 41 ] ? r - ( 60'd1 << 54 ) : r ;
         r = b [ 40 ] ? r - ( 60'd1 << 53 ) : r ;
         r = b [ 39 ] ? r - ( 60'd1 << 52 ) : r ;
         r = b [ 38 ] ? r - ( 60'd1 << 51 ) : r ;
         r = b [ 37 ] ? r - ( 60'd1 << 50 ) : r ;
         r = b [ 36 ] ? r - ( 60'd1 << 49 ) : r ;
         r = b [ 35 ] ? r - ( 60'd1 << 48 ) : r ;
         r = b [ 34 ] ? r - ( 60'd1 << 47 ) : r ;
         r = b [ 33 ] ? r - ( 60'd1 << 46 ) : r ;
         r = b [ 32 ] ? r - ( 60'd1 << 45 ) : r ;
         r = b [ 31 ] ? r - ( 60'd1 << 44 ) : r ;
         r = b [ 30 ] ? r - ( 60'd1 << 43 ) : r ;
         r = b [ 29 ] ? r - ( 60'd1 << 42 ) : r ;
         r = b [ 28 ] ? r - ( 60'd1 << 41 ) : r ;
         r = b [ 27 ] ? r - ( 60'd1 << 40 ) : r ;
         r = b [ 26 ] ? r - ( 60'd1 << 39 ) : r ;
         r = b [ 25 ] ? r - ( 60'd1 << 38 ) : r ;
         r = b [ 24 ] ? r - ( 60'd1 << 37 ) : r ;
         r = b [ 23 ] ? r - ( 60'd1 << 36 ) : r ;
         r = b [ 22 ] ? r - ( 60'd1 << 35 ) : r ;
         r = b [ 21 ] ? r - ( 60'd1 << 34 ) : r ;
         r = b [ 20 ] ? r - ( 60'd1 << 33 ) : r ;
         r = b [ 19 ] ? r - ( 60'd1 << 32 ) : r ;
         r = b [ 18 ] ? r - ( 60'd1 << 31 ) : r ;
         r = b [ 17 ] ? r - ( 60'd1 << 30 ) : r ;
         r = b [ 16 ] ? r - ( 60'd1 << 29 ) : r ;
         r = b [ 15 ] ? r - ( 60'd1 << 28 ) : r ;
         r = b [ 14 ] ? r - ( 60'd1 << 27 ) : r ;
         r = b [ 13 ] ? r - ( 60'd1 << 26 ) : r ;
         r = b [ 12 ] ? r - ( 60'd1 << 25 ) : r ;
         r = b [ 11 ] ? r - ( 60'd1 << 24 ) : r ;
         r = b [ 10 ] ? r - ( 60'd1 << 23 ) : r ;
         r = b [ 9 ] ? r - ( 60'd1 << 22 ) : r ;
         r = b [ 8 ] ? r - ( 60'd1 << 21 ) : r ;
         r = b [ 7 ] ? r - ( 60'd1 << 20 ) : r ;
         r = b [ 6 ] ? r - ( 60'd1 << 19 ) : r ;
         r = b [ 5 ] ? r - ( 60'd1 << 18 ) : r ;
         r = b [ 4 ] ? r - ( 60'd1 << 17 ) : r ;
         r = b [ 3 ] ? r - ( 60'd1 << 16 ) : r ;
         r = b [ 2 ] ? r - ( 60'd1 << 15 ) : r ;
         r = b [ 1 ] ? r - ( 60'd1 << 14 ) : r ;
         r = b [ 0 ] ? r - ( 60'd1 << 13 ) : r ;
      end

// Bit by Bit Multiply & Divide + Modulus
// Copyright © 2022 by Gregory Scott Callen
// All Rights Reserved.

      if (( b << 12n ) <= r ) begin
         n = n | 60'd4096;
         r = b [ 47 ] ? r - ( 60'd1 << 59 ) : r ;
         r = b [ 46 ] ? r - ( 60'd1 << 58 ) : r ;
         r = b [ 45 ] ? r - ( 60'd1 << 57 ) : r ;
         r = b [ 44 ] ? r - ( 60'd1 << 56 ) : r ;
         r = b [ 43 ] ? r - ( 60'd1 << 55 ) : r ;
         r = b [ 42 ] ? r - ( 60'd1 << 54 ) : r ;
         r = b [ 41 ] ? r - ( 60'd1 << 53 ) : r ;
         r = b [ 40 ] ? r - ( 60'd1 << 52 ) : r ;
         r = b [ 39 ] ? r - ( 60'd1 << 51 ) : r ;
         r = b [ 38 ] ? r - ( 60'd1 << 50 ) : r ;
         r = b [ 37 ] ? r - ( 60'd1 << 49 ) : r ;
         r = b [ 36 ] ? r - ( 60'd1 << 48 ) : r ;
         r = b [ 35 ] ? r - ( 60'd1 << 47 ) : r ;
         r = b [ 34 ] ? r - ( 60'd1 << 46 ) : r ;
         r = b [ 33 ] ? r - ( 60'd1 << 45 ) : r ;
         r = b [ 32 ] ? r - ( 60'd1 << 44 ) : r ;
         r = b [ 31 ] ? r - ( 60'd1 << 43 ) : r ;
         r = b [ 30 ] ? r - ( 60'd1 << 42 ) : r ;
         r = b [ 29 ] ? r - ( 60'd1 << 41 ) : r ;
         r = b [ 28 ] ? r - ( 60'd1 << 40 ) : r ;
         r = b [ 27 ] ? r - ( 60'd1 << 39 ) : r ;
         r = b [ 26 ] ? r - ( 60'd1 << 38 ) : r ;
         r = b [ 25 ] ? r - ( 60'd1 << 37 ) : r ;
         r = b [ 24 ] ? r - ( 60'd1 << 36 ) : r ;
         r = b [ 23 ] ? r - ( 60'd1 << 35 ) : r ;
         r = b [ 22 ] ? r - ( 60'd1 << 34 ) : r ;
         r = b [ 21 ] ? r - ( 60'd1 << 33 ) : r ;
         r = b [ 20 ] ? r - ( 60'd1 << 32 ) : r ;
         r = b [ 19 ] ? r - ( 60'd1 << 31 ) : r ;
         r = b [ 18 ] ? r - ( 60'd1 << 30 ) : r ;
         r = b [ 17 ] ? r - ( 60'd1 << 29 ) : r ;
         r = b [ 16 ] ? r - ( 60'd1 << 28 ) : r ;
         r = b [ 15 ] ? r - ( 60'd1 << 27 ) : r ;
         r = b [ 14 ] ? r - ( 60'd1 << 26 ) : r ;
         r = b [ 13 ] ? r - ( 60'd1 << 25 ) : r ;
         r = b [ 12 ] ? r - ( 60'd1 << 24 ) : r ;
         r = b [ 11 ] ? r - ( 60'd1 << 23 ) : r ;
         r = b [ 10 ] ? r - ( 60'd1 << 22 ) : r ;
         r = b [ 9 ] ? r - ( 60'd1 << 21 ) : r ;
         r = b [ 8 ] ? r - ( 60'd1 << 20 ) : r ;
         r = b [ 7 ] ? r - ( 60'd1 << 19 ) : r ;
         r = b [ 6 ] ? r - ( 60'd1 << 18 ) : r ;
         r = b [ 5 ] ? r - ( 60'd1 << 17 ) : r ;
         r = b [ 4 ] ? r - ( 60'd1 << 16 ) : r ;
         r = b [ 3 ] ? r - ( 60'd1 << 15 ) : r ;
         r = b [ 2 ] ? r - ( 60'd1 << 14 ) : r ;
         r = b [ 1 ] ? r - ( 60'd1 << 13 ) : r ;
         r = b [ 0 ] ? r - ( 60'd1 << 12 ) : r ;
      end

// Bit by Bit Multiply & Divide + Modulus
// Copyright © 2022 by Gregory Scott Callen
// All Rights Reserved.

      if (( b << 11n ) <= r ) begin
         n = n | 60'd2048;
         r = b [ 48 ] ? r - ( 60'd1 << 59 ) : r ;
         r = b [ 47 ] ? r - ( 60'd1 << 58 ) : r ;
         r = b [ 46 ] ? r - ( 60'd1 << 57 ) : r ;
         r = b [ 45 ] ? r - ( 60'd1 << 56 ) : r ;
         r = b [ 44 ] ? r - ( 60'd1 << 55 ) : r ;
         r = b [ 43 ] ? r - ( 60'd1 << 54 ) : r ;
         r = b [ 42 ] ? r - ( 60'd1 << 53 ) : r ;
         r = b [ 41 ] ? r - ( 60'd1 << 52 ) : r ;
         r = b [ 40 ] ? r - ( 60'd1 << 51 ) : r ;
         r = b [ 39 ] ? r - ( 60'd1 << 50 ) : r ;
         r = b [ 38 ] ? r - ( 60'd1 << 49 ) : r ;
         r = b [ 37 ] ? r - ( 60'd1 << 48 ) : r ;
         r = b [ 36 ] ? r - ( 60'd1 << 47 ) : r ;
         r = b [ 35 ] ? r - ( 60'd1 << 46 ) : r ;
         r = b [ 34 ] ? r - ( 60'd1 << 45 ) : r ;
         r = b [ 33 ] ? r - ( 60'd1 << 44 ) : r ;
         r = b [ 32 ] ? r - ( 60'd1 << 43 ) : r ;
         r = b [ 31 ] ? r - ( 60'd1 << 42 ) : r ;
         r = b [ 30 ] ? r - ( 60'd1 << 41 ) : r ;
         r = b [ 29 ] ? r - ( 60'd1 << 40 ) : r ;
         r = b [ 28 ] ? r - ( 60'd1 << 39 ) : r ;
         r = b [ 27 ] ? r - ( 60'd1 << 38 ) : r ;
         r = b [ 26 ] ? r - ( 60'd1 << 37 ) : r ;
         r = b [ 25 ] ? r - ( 60'd1 << 36 ) : r ;
         r = b [ 24 ] ? r - ( 60'd1 << 35 ) : r ;
         r = b [ 23 ] ? r - ( 60'd1 << 34 ) : r ;
         r = b [ 22 ] ? r - ( 60'd1 << 33 ) : r ;
         r = b [ 21 ] ? r - ( 60'd1 << 32 ) : r ;
         r = b [ 20 ] ? r - ( 60'd1 << 31 ) : r ;
         r = b [ 19 ] ? r - ( 60'd1 << 30 ) : r ;
         r = b [ 18 ] ? r - ( 60'd1 << 29 ) : r ;
         r = b [ 17 ] ? r - ( 60'd1 << 28 ) : r ;
         r = b [ 16 ] ? r - ( 60'd1 << 27 ) : r ;
         r = b [ 15 ] ? r - ( 60'd1 << 26 ) : r ;
         r = b [ 14 ] ? r - ( 60'd1 << 25 ) : r ;
         r = b [ 13 ] ? r - ( 60'd1 << 24 ) : r ;
         r = b [ 12 ] ? r - ( 60'd1 << 23 ) : r ;
         r = b [ 11 ] ? r - ( 60'd1 << 22 ) : r ;
         r = b [ 10 ] ? r - ( 60'd1 << 21 ) : r ;
         r = b [ 9 ] ? r - ( 60'd1 << 20 ) : r ;
         r = b [ 8 ] ? r - ( 60'd1 << 19 ) : r ;
         r = b [ 7 ] ? r - ( 60'd1 << 18 ) : r ;
         r = b [ 6 ] ? r - ( 60'd1 << 17 ) : r ;
         r = b [ 5 ] ? r - ( 60'd1 << 16 ) : r ;
         r = b [ 4 ] ? r - ( 60'd1 << 15 ) : r ;
         r = b [ 3 ] ? r - ( 60'd1 << 14 ) : r ;
         r = b [ 2 ] ? r - ( 60'd1 << 13 ) : r ;
         r = b [ 1 ] ? r - ( 60'd1 << 12 ) : r ;
         r = b [ 0 ] ? r - ( 60'd1 << 11 ) : r ;
      end

// Bit by Bit Multiply & Divide + Modulus
// Copyright © 2022 by Gregory Scott Callen
// All Rights Reserved.

      if (( b << 10n ) <= r ) begin
         n = n | 60'd1024;
         r = b [ 49 ] ? r - ( 60'd1 << 59 ) : r ;
         r = b [ 48 ] ? r - ( 60'd1 << 58 ) : r ;
         r = b [ 47 ] ? r - ( 60'd1 << 57 ) : r ;
         r = b [ 46 ] ? r - ( 60'd1 << 56 ) : r ;
         r = b [ 45 ] ? r - ( 60'd1 << 55 ) : r ;
         r = b [ 44 ] ? r - ( 60'd1 << 54 ) : r ;
         r = b [ 43 ] ? r - ( 60'd1 << 53 ) : r ;
         r = b [ 42 ] ? r - ( 60'd1 << 52 ) : r ;
         r = b [ 41 ] ? r - ( 60'd1 << 51 ) : r ;
         r = b [ 40 ] ? r - ( 60'd1 << 50 ) : r ;
         r = b [ 39 ] ? r - ( 60'd1 << 49 ) : r ;
         r = b [ 38 ] ? r - ( 60'd1 << 48 ) : r ;
         r = b [ 37 ] ? r - ( 60'd1 << 47 ) : r ;
         r = b [ 36 ] ? r - ( 60'd1 << 46 ) : r ;
         r = b [ 35 ] ? r - ( 60'd1 << 45 ) : r ;
         r = b [ 34 ] ? r - ( 60'd1 << 44 ) : r ;
         r = b [ 33 ] ? r - ( 60'd1 << 43 ) : r ;
         r = b [ 32 ] ? r - ( 60'd1 << 42 ) : r ;
         r = b [ 31 ] ? r - ( 60'd1 << 41 ) : r ;
         r = b [ 30 ] ? r - ( 60'd1 << 40 ) : r ;
         r = b [ 29 ] ? r - ( 60'd1 << 39 ) : r ;
         r = b [ 28 ] ? r - ( 60'd1 << 38 ) : r ;
         r = b [ 27 ] ? r - ( 60'd1 << 37 ) : r ;
         r = b [ 26 ] ? r - ( 60'd1 << 36 ) : r ;
         r = b [ 25 ] ? r - ( 60'd1 << 35 ) : r ;
         r = b [ 24 ] ? r - ( 60'd1 << 34 ) : r ;
         r = b [ 23 ] ? r - ( 60'd1 << 33 ) : r ;
         r = b [ 22 ] ? r - ( 60'd1 << 32 ) : r ;
         r = b [ 21 ] ? r - ( 60'd1 << 31 ) : r ;
         r = b [ 20 ] ? r - ( 60'd1 << 30 ) : r ;
         r = b [ 19 ] ? r - ( 60'd1 << 29 ) : r ;
         r = b [ 18 ] ? r - ( 60'd1 << 28 ) : r ;
         r = b [ 17 ] ? r - ( 60'd1 << 27 ) : r ;
         r = b [ 16 ] ? r - ( 60'd1 << 26 ) : r ;
         r = b [ 15 ] ? r - ( 60'd1 << 25 ) : r ;
         r = b [ 14 ] ? r - ( 60'd1 << 24 ) : r ;
         r = b [ 13 ] ? r - ( 60'd1 << 23 ) : r ;
         r = b [ 12 ] ? r - ( 60'd1 << 22 ) : r ;
         r = b [ 11 ] ? r - ( 60'd1 << 21 ) : r ;
         r = b [ 10 ] ? r - ( 60'd1 << 20 ) : r ;
         r = b [ 9 ] ? r - ( 60'd1 << 19 ) : r ;
         r = b [ 8 ] ? r - ( 60'd1 << 18 ) : r ;
         r = b [ 7 ] ? r - ( 60'd1 << 17 ) : r ;
         r = b [ 6 ] ? r - ( 60'd1 << 16 ) : r ;
         r = b [ 5 ] ? r - ( 60'd1 << 15 ) : r ;
         r = b [ 4 ] ? r - ( 60'd1 << 14 ) : r ;
         r = b [ 3 ] ? r - ( 60'd1 << 13 ) : r ;
         r = b [ 2 ] ? r - ( 60'd1 << 12 ) : r ;
         r = b [ 1 ] ? r - ( 60'd1 << 11 ) : r ;
         r = b [ 0 ] ? r - ( 60'd1 << 10 ) : r ;
      end

// Bit by Bit Multiply & Divide + Modulus
// Copyright © 2022 by Gregory Scott Callen
// All Rights Reserved.

      if (( b << 9n ) <= r ) begin
         n = n | 60'd512;
         r = b [ 50 ] ? r - ( 60'd1 << 59 ) : r ;
         r = b [ 49 ] ? r - ( 60'd1 << 58 ) : r ;
         r = b [ 48 ] ? r - ( 60'd1 << 57 ) : r ;
         r = b [ 47 ] ? r - ( 60'd1 << 56 ) : r ;
         r = b [ 46 ] ? r - ( 60'd1 << 55 ) : r ;
         r = b [ 45 ] ? r - ( 60'd1 << 54 ) : r ;
         r = b [ 44 ] ? r - ( 60'd1 << 53 ) : r ;
         r = b [ 43 ] ? r - ( 60'd1 << 52 ) : r ;
         r = b [ 42 ] ? r - ( 60'd1 << 51 ) : r ;
         r = b [ 41 ] ? r - ( 60'd1 << 50 ) : r ;
         r = b [ 40 ] ? r - ( 60'd1 << 49 ) : r ;
         r = b [ 39 ] ? r - ( 60'd1 << 48 ) : r ;
         r = b [ 38 ] ? r - ( 60'd1 << 47 ) : r ;
         r = b [ 37 ] ? r - ( 60'd1 << 46 ) : r ;
         r = b [ 36 ] ? r - ( 60'd1 << 45 ) : r ;
         r = b [ 35 ] ? r - ( 60'd1 << 44 ) : r ;
         r = b [ 34 ] ? r - ( 60'd1 << 43 ) : r ;
         r = b [ 33 ] ? r - ( 60'd1 << 42 ) : r ;
         r = b [ 32 ] ? r - ( 60'd1 << 41 ) : r ;
         r = b [ 31 ] ? r - ( 60'd1 << 40 ) : r ;
         r = b [ 30 ] ? r - ( 60'd1 << 39 ) : r ;
         r = b [ 29 ] ? r - ( 60'd1 << 38 ) : r ;
         r = b [ 28 ] ? r - ( 60'd1 << 37 ) : r ;
         r = b [ 27 ] ? r - ( 60'd1 << 36 ) : r ;
         r = b [ 26 ] ? r - ( 60'd1 << 35 ) : r ;
         r = b [ 25 ] ? r - ( 60'd1 << 34 ) : r ;
         r = b [ 24 ] ? r - ( 60'd1 << 33 ) : r ;
         r = b [ 23 ] ? r - ( 60'd1 << 32 ) : r ;
         r = b [ 22 ] ? r - ( 60'd1 << 31 ) : r ;
         r = b [ 21 ] ? r - ( 60'd1 << 30 ) : r ;
         r = b [ 20 ] ? r - ( 60'd1 << 29 ) : r ;
         r = b [ 19 ] ? r - ( 60'd1 << 28 ) : r ;
         r = b [ 18 ] ? r - ( 60'd1 << 27 ) : r ;
         r = b [ 17 ] ? r - ( 60'd1 << 26 ) : r ;
         r = b [ 16 ] ? r - ( 60'd1 << 25 ) : r ;
         r = b [ 15 ] ? r - ( 60'd1 << 24 ) : r ;
         r = b [ 14 ] ? r - ( 60'd1 << 23 ) : r ;
         r = b [ 13 ] ? r - ( 60'd1 << 22 ) : r ;
         r = b [ 12 ] ? r - ( 60'd1 << 21 ) : r ;
         r = b [ 11 ] ? r - ( 60'd1 << 20 ) : r ;
         r = b [ 10 ] ? r - ( 60'd1 << 19 ) : r ;
         r = b [ 9 ] ? r - ( 60'd1 << 18 ) : r ;
         r = b [ 8 ] ? r - ( 60'd1 << 17 ) : r ;
         r = b [ 7 ] ? r - ( 60'd1 << 16 ) : r ;
         r = b [ 6 ] ? r - ( 60'd1 << 15 ) : r ;
         r = b [ 5 ] ? r - ( 60'd1 << 14 ) : r ;
         r = b [ 4 ] ? r - ( 60'd1 << 13 ) : r ;
         r = b [ 3 ] ? r - ( 60'd1 << 12 ) : r ;
         r = b [ 2 ] ? r - ( 60'd1 << 11 ) : r ;
         r = b [ 1 ] ? r - ( 60'd1 << 10 ) : r ;
         r = b [ 0 ] ? r - ( 60'd1 << 9 ) : r ;
      end

// Bit by Bit Multiply & Divide + Modulus
// Copyright © 2022 by Gregory Scott Callen
// All Rights Reserved.

      if (( b << 8n ) <= r ) begin
         n = n | 60'd256;
         r = b [ 51 ] ? r - ( 60'd1 << 59 ) : r ;
         r = b [ 50 ] ? r - ( 60'd1 << 58 ) : r ;
         r = b [ 49 ] ? r - ( 60'd1 << 57 ) : r ;
         r = b [ 48 ] ? r - ( 60'd1 << 56 ) : r ;
         r = b [ 47 ] ? r - ( 60'd1 << 55 ) : r ;
         r = b [ 46 ] ? r - ( 60'd1 << 54 ) : r ;
         r = b [ 45 ] ? r - ( 60'd1 << 53 ) : r ;
         r = b [ 44 ] ? r - ( 60'd1 << 52 ) : r ;
         r = b [ 43 ] ? r - ( 60'd1 << 51 ) : r ;
         r = b [ 42 ] ? r - ( 60'd1 << 50 ) : r ;
         r = b [ 41 ] ? r - ( 60'd1 << 49 ) : r ;
         r = b [ 40 ] ? r - ( 60'd1 << 48 ) : r ;
         r = b [ 39 ] ? r - ( 60'd1 << 47 ) : r ;
         r = b [ 38 ] ? r - ( 60'd1 << 46 ) : r ;
         r = b [ 37 ] ? r - ( 60'd1 << 45 ) : r ;
         r = b [ 36 ] ? r - ( 60'd1 << 44 ) : r ;
         r = b [ 35 ] ? r - ( 60'd1 << 43 ) : r ;
         r = b [ 34 ] ? r - ( 60'd1 << 42 ) : r ;
         r = b [ 33 ] ? r - ( 60'd1 << 41 ) : r ;
         r = b [ 32 ] ? r - ( 60'd1 << 40 ) : r ;
         r = b [ 31 ] ? r - ( 60'd1 << 39 ) : r ;
         r = b [ 30 ] ? r - ( 60'd1 << 38 ) : r ;
         r = b [ 29 ] ? r - ( 60'd1 << 37 ) : r ;
         r = b [ 28 ] ? r - ( 60'd1 << 36 ) : r ;
         r = b [ 27 ] ? r - ( 60'd1 << 35 ) : r ;
         r = b [ 26 ] ? r - ( 60'd1 << 34 ) : r ;
         r = b [ 25 ] ? r - ( 60'd1 << 33 ) : r ;
         r = b [ 24 ] ? r - ( 60'd1 << 32 ) : r ;
         r = b [ 23 ] ? r - ( 60'd1 << 31 ) : r ;
         r = b [ 22 ] ? r - ( 60'd1 << 30 ) : r ;
         r = b [ 21 ] ? r - ( 60'd1 << 29 ) : r ;
         r = b [ 20 ] ? r - ( 60'd1 << 28 ) : r ;
         r = b [ 19 ] ? r - ( 60'd1 << 27 ) : r ;
         r = b [ 18 ] ? r - ( 60'd1 << 26 ) : r ;
         r = b [ 17 ] ? r - ( 60'd1 << 25 ) : r ;
         r = b [ 16 ] ? r - ( 60'd1 << 24 ) : r ;
         r = b [ 15 ] ? r - ( 60'd1 << 23 ) : r ;
         r = b [ 14 ] ? r - ( 60'd1 << 22 ) : r ;
         r = b [ 13 ] ? r - ( 60'd1 << 21 ) : r ;
         r = b [ 12 ] ? r - ( 60'd1 << 20 ) : r ;
         r = b [ 11 ] ? r - ( 60'd1 << 19 ) : r ;
         r = b [ 10 ] ? r - ( 60'd1 << 18 ) : r ;
         r = b [ 9 ] ? r - ( 60'd1 << 17 ) : r ;
         r = b [ 8 ] ? r - ( 60'd1 << 16 ) : r ;
         r = b [ 7 ] ? r - ( 60'd1 << 15 ) : r ;
         r = b [ 6 ] ? r - ( 60'd1 << 14 ) : r ;
         r = b [ 5 ] ? r - ( 60'd1 << 13 ) : r ;
         r = b [ 4 ] ? r - ( 60'd1 << 12 ) : r ;
         r = b [ 3 ] ? r - ( 60'd1 << 11 ) : r ;
         r = b [ 2 ] ? r - ( 60'd1 << 10 ) : r ;
         r = b [ 1 ] ? r - ( 60'd1 << 9 ) : r ;
         r = b [ 0 ] ? r - ( 60'd1 << 8 ) : r ;
      end

// Bit by Bit Multiply & Divide + Modulus
// Copyright © 2022 by Gregory Scott Callen
// All Rights Reserved.

      if (( b << 7n ) <= r ) begin
         n = n | 60'd128;
         r = b [ 52 ] ? r - ( 60'd1 << 59 ) : r ;
         r = b [ 51 ] ? r - ( 60'd1 << 58 ) : r ;
         r = b [ 50 ] ? r - ( 60'd1 << 57 ) : r ;
         r = b [ 49 ] ? r - ( 60'd1 << 56 ) : r ;
         r = b [ 48 ] ? r - ( 60'd1 << 55 ) : r ;
         r = b [ 47 ] ? r - ( 60'd1 << 54 ) : r ;
         r = b [ 46 ] ? r - ( 60'd1 << 53 ) : r ;
         r = b [ 45 ] ? r - ( 60'd1 << 52 ) : r ;
         r = b [ 44 ] ? r - ( 60'd1 << 51 ) : r ;
         r = b [ 43 ] ? r - ( 60'd1 << 50 ) : r ;
         r = b [ 42 ] ? r - ( 60'd1 << 49 ) : r ;
         r = b [ 41 ] ? r - ( 60'd1 << 48 ) : r ;
         r = b [ 40 ] ? r - ( 60'd1 << 47 ) : r ;
         r = b [ 39 ] ? r - ( 60'd1 << 46 ) : r ;
         r = b [ 38 ] ? r - ( 60'd1 << 45 ) : r ;
         r = b [ 37 ] ? r - ( 60'd1 << 44 ) : r ;
         r = b [ 36 ] ? r - ( 60'd1 << 43 ) : r ;
         r = b [ 35 ] ? r - ( 60'd1 << 42 ) : r ;
         r = b [ 34 ] ? r - ( 60'd1 << 41 ) : r ;
         r = b [ 33 ] ? r - ( 60'd1 << 40 ) : r ;
         r = b [ 32 ] ? r - ( 60'd1 << 39 ) : r ;
         r = b [ 31 ] ? r - ( 60'd1 << 38 ) : r ;
         r = b [ 30 ] ? r - ( 60'd1 << 37 ) : r ;
         r = b [ 29 ] ? r - ( 60'd1 << 36 ) : r ;
         r = b [ 28 ] ? r - ( 60'd1 << 35 ) : r ;
         r = b [ 27 ] ? r - ( 60'd1 << 34 ) : r ;
         r = b [ 26 ] ? r - ( 60'd1 << 33 ) : r ;
         r = b [ 25 ] ? r - ( 60'd1 << 32 ) : r ;
         r = b [ 24 ] ? r - ( 60'd1 << 31 ) : r ;
         r = b [ 23 ] ? r - ( 60'd1 << 30 ) : r ;
         r = b [ 22 ] ? r - ( 60'd1 << 29 ) : r ;
         r = b [ 21 ] ? r - ( 60'd1 << 28 ) : r ;
         r = b [ 20 ] ? r - ( 60'd1 << 27 ) : r ;
         r = b [ 19 ] ? r - ( 60'd1 << 26 ) : r ;
         r = b [ 18 ] ? r - ( 60'd1 << 25 ) : r ;
         r = b [ 17 ] ? r - ( 60'd1 << 24 ) : r ;
         r = b [ 16 ] ? r - ( 60'd1 << 23 ) : r ;
         r = b [ 15 ] ? r - ( 60'd1 << 22 ) : r ;
         r = b [ 14 ] ? r - ( 60'd1 << 21 ) : r ;
         r = b [ 13 ] ? r - ( 60'd1 << 20 ) : r ;
         r = b [ 12 ] ? r - ( 60'd1 << 19 ) : r ;
         r = b [ 11 ] ? r - ( 60'd1 << 18 ) : r ;
         r = b [ 10 ] ? r - ( 60'd1 << 17 ) : r ;
         r = b [ 9 ] ? r - ( 60'd1 << 16 ) : r ;
         r = b [ 8 ] ? r - ( 60'd1 << 15 ) : r ;
         r = b [ 7 ] ? r - ( 60'd1 << 14 ) : r ;
         r = b [ 6 ] ? r - ( 60'd1 << 13 ) : r ;
         r = b [ 5 ] ? r - ( 60'd1 << 12 ) : r ;
         r = b [ 4 ] ? r - ( 60'd1 << 11 ) : r ;
         r = b [ 3 ] ? r - ( 60'd1 << 10 ) : r ;
         r = b [ 2 ] ? r - ( 60'd1 << 9 ) : r ;
         r = b [ 1 ] ? r - ( 60'd1 << 8 ) : r ;
         r = b [ 0 ] ? r - ( 60'd1 << 7 ) : r ;
      end

// Bit by Bit Multiply & Divide + Modulus
// Copyright © 2022 by Gregory Scott Callen
// All Rights Reserved.

      if (( b << 6n ) <= r ) begin
         n = n | 60'd64;
         r = b [ 53 ] ? r - ( 60'd1 << 59 ) : r ;
         r = b [ 52 ] ? r - ( 60'd1 << 58 ) : r ;
         r = b [ 51 ] ? r - ( 60'd1 << 57 ) : r ;
         r = b [ 50 ] ? r - ( 60'd1 << 56 ) : r ;
         r = b [ 49 ] ? r - ( 60'd1 << 55 ) : r ;
         r = b [ 48 ] ? r - ( 60'd1 << 54 ) : r ;
         r = b [ 47 ] ? r - ( 60'd1 << 53 ) : r ;
         r = b [ 46 ] ? r - ( 60'd1 << 52 ) : r ;
         r = b [ 45 ] ? r - ( 60'd1 << 51 ) : r ;
         r = b [ 44 ] ? r - ( 60'd1 << 50 ) : r ;
         r = b [ 43 ] ? r - ( 60'd1 << 49 ) : r ;
         r = b [ 42 ] ? r - ( 60'd1 << 48 ) : r ;
         r = b [ 41 ] ? r - ( 60'd1 << 47 ) : r ;
         r = b [ 40 ] ? r - ( 60'd1 << 46 ) : r ;
         r = b [ 39 ] ? r - ( 60'd1 << 45 ) : r ;
         r = b [ 38 ] ? r - ( 60'd1 << 44 ) : r ;
         r = b [ 37 ] ? r - ( 60'd1 << 43 ) : r ;
         r = b [ 36 ] ? r - ( 60'd1 << 42 ) : r ;
         r = b [ 35 ] ? r - ( 60'd1 << 41 ) : r ;
         r = b [ 34 ] ? r - ( 60'd1 << 40 ) : r ;
         r = b [ 33 ] ? r - ( 60'd1 << 39 ) : r ;
         r = b [ 32 ] ? r - ( 60'd1 << 38 ) : r ;
         r = b [ 31 ] ? r - ( 60'd1 << 37 ) : r ;
         r = b [ 30 ] ? r - ( 60'd1 << 36 ) : r ;
         r = b [ 29 ] ? r - ( 60'd1 << 35 ) : r ;
         r = b [ 28 ] ? r - ( 60'd1 << 34 ) : r ;
         r = b [ 27 ] ? r - ( 60'd1 << 33 ) : r ;
         r = b [ 26 ] ? r - ( 60'd1 << 32 ) : r ;
         r = b [ 25 ] ? r - ( 60'd1 << 31 ) : r ;
         r = b [ 24 ] ? r - ( 60'd1 << 30 ) : r ;
         r = b [ 23 ] ? r - ( 60'd1 << 29 ) : r ;
         r = b [ 22 ] ? r - ( 60'd1 << 28 ) : r ;
         r = b [ 21 ] ? r - ( 60'd1 << 27 ) : r ;
         r = b [ 20 ] ? r - ( 60'd1 << 26 ) : r ;
         r = b [ 19 ] ? r - ( 60'd1 << 25 ) : r ;
         r = b [ 18 ] ? r - ( 60'd1 << 24 ) : r ;
         r = b [ 17 ] ? r - ( 60'd1 << 23 ) : r ;
         r = b [ 16 ] ? r - ( 60'd1 << 22 ) : r ;
         r = b [ 15 ] ? r - ( 60'd1 << 21 ) : r ;
         r = b [ 14 ] ? r - ( 60'd1 << 20 ) : r ;
         r = b [ 13 ] ? r - ( 60'd1 << 19 ) : r ;
         r = b [ 12 ] ? r - ( 60'd1 << 18 ) : r ;
         r = b [ 11 ] ? r - ( 60'd1 << 17 ) : r ;
         r = b [ 10 ] ? r - ( 60'd1 << 16 ) : r ;
         r = b [ 9 ] ? r - ( 60'd1 << 15 ) : r ;
         r = b [ 8 ] ? r - ( 60'd1 << 14 ) : r ;
         r = b [ 7 ] ? r - ( 60'd1 << 13 ) : r ;
         r = b [ 6 ] ? r - ( 60'd1 << 12 ) : r ;
         r = b [ 5 ] ? r - ( 60'd1 << 11 ) : r ;
         r = b [ 4 ] ? r - ( 60'd1 << 10 ) : r ;
         r = b [ 3 ] ? r - ( 60'd1 << 9 ) : r ;
         r = b [ 2 ] ? r - ( 60'd1 << 8 ) : r ;
         r = b [ 1 ] ? r - ( 60'd1 << 7 ) : r ;
         r = b [ 0 ] ? r - ( 60'd1 << 6 ) : r ;
      end

// Bit by Bit Multiply & Divide + Modulus
// Copyright © 2022 by Gregory Scott Callen
// All Rights Reserved.

      if (( b << 5n ) <= r ) begin
         n = n | 60'd32;
         r = b [ 54 ] ? r - ( 60'd1 << 59 ) : r ;
         r = b [ 53 ] ? r - ( 60'd1 << 58 ) : r ;
         r = b [ 52 ] ? r - ( 60'd1 << 57 ) : r ;
         r = b [ 51 ] ? r - ( 60'd1 << 56 ) : r ;
         r = b [ 50 ] ? r - ( 60'd1 << 55 ) : r ;
         r = b [ 49 ] ? r - ( 60'd1 << 54 ) : r ;
         r = b [ 48 ] ? r - ( 60'd1 << 53 ) : r ;
         r = b [ 47 ] ? r - ( 60'd1 << 52 ) : r ;
         r = b [ 46 ] ? r - ( 60'd1 << 51 ) : r ;
         r = b [ 45 ] ? r - ( 60'd1 << 50 ) : r ;
         r = b [ 44 ] ? r - ( 60'd1 << 49 ) : r ;
         r = b [ 43 ] ? r - ( 60'd1 << 48 ) : r ;
         r = b [ 42 ] ? r - ( 60'd1 << 47 ) : r ;
         r = b [ 41 ] ? r - ( 60'd1 << 46 ) : r ;
         r = b [ 40 ] ? r - ( 60'd1 << 45 ) : r ;
         r = b [ 39 ] ? r - ( 60'd1 << 44 ) : r ;
         r = b [ 38 ] ? r - ( 60'd1 << 43 ) : r ;
         r = b [ 37 ] ? r - ( 60'd1 << 42 ) : r ;
         r = b [ 36 ] ? r - ( 60'd1 << 41 ) : r ;
         r = b [ 35 ] ? r - ( 60'd1 << 40 ) : r ;
         r = b [ 34 ] ? r - ( 60'd1 << 39 ) : r ;
         r = b [ 33 ] ? r - ( 60'd1 << 38 ) : r ;
         r = b [ 32 ] ? r - ( 60'd1 << 37 ) : r ;
         r = b [ 31 ] ? r - ( 60'd1 << 36 ) : r ;
         r = b [ 30 ] ? r - ( 60'd1 << 35 ) : r ;
         r = b [ 29 ] ? r - ( 60'd1 << 34 ) : r ;
         r = b [ 28 ] ? r - ( 60'd1 << 33 ) : r ;
         r = b [ 27 ] ? r - ( 60'd1 << 32 ) : r ;
         r = b [ 26 ] ? r - ( 60'd1 << 31 ) : r ;
         r = b [ 25 ] ? r - ( 60'd1 << 30 ) : r ;
         r = b [ 24 ] ? r - ( 60'd1 << 29 ) : r ;
         r = b [ 23 ] ? r - ( 60'd1 << 28 ) : r ;
         r = b [ 22 ] ? r - ( 60'd1 << 27 ) : r ;
         r = b [ 21 ] ? r - ( 60'd1 << 26 ) : r ;
         r = b [ 20 ] ? r - ( 60'd1 << 25 ) : r ;
         r = b [ 19 ] ? r - ( 60'd1 << 24 ) : r ;
         r = b [ 18 ] ? r - ( 60'd1 << 23 ) : r ;
         r = b [ 17 ] ? r - ( 60'd1 << 22 ) : r ;
         r = b [ 16 ] ? r - ( 60'd1 << 21 ) : r ;
         r = b [ 15 ] ? r - ( 60'd1 << 20 ) : r ;
         r = b [ 14 ] ? r - ( 60'd1 << 19 ) : r ;
         r = b [ 13 ] ? r - ( 60'd1 << 18 ) : r ;
         r = b [ 12 ] ? r - ( 60'd1 << 17 ) : r ;
         r = b [ 11 ] ? r - ( 60'd1 << 16 ) : r ;
         r = b [ 10 ] ? r - ( 60'd1 << 15 ) : r ;
         r = b [ 9 ] ? r - ( 60'd1 << 14 ) : r ;
         r = b [ 8 ] ? r - ( 60'd1 << 13 ) : r ;
         r = b [ 7 ] ? r - ( 60'd1 << 12 ) : r ;
         r = b [ 6 ] ? r - ( 60'd1 << 11 ) : r ;
         r = b [ 5 ] ? r - ( 60'd1 << 10 ) : r ;
         r = b [ 4 ] ? r - ( 60'd1 << 9 ) : r ;
         r = b [ 3 ] ? r - ( 60'd1 << 8 ) : r ;
         r = b [ 2 ] ? r - ( 60'd1 << 7 ) : r ;
         r = b [ 1 ] ? r - ( 60'd1 << 6 ) : r ;
         r = b [ 0 ] ? r - ( 60'd1 << 5 ) : r ;
      end

// Bit by Bit Multiply & Divide + Modulus
// Copyright © 2022 by Gregory Scott Callen
// All Rights Reserved.

      if (( b << 4n ) <= r ) begin
         n = n | 60'd16;
         r = b [ 55 ] ? r - ( 60'd1 << 59 ) : r ;
         r = b [ 54 ] ? r - ( 60'd1 << 58 ) : r ;
         r = b [ 53 ] ? r - ( 60'd1 << 57 ) : r ;
         r = b [ 52 ] ? r - ( 60'd1 << 56 ) : r ;
         r = b [ 51 ] ? r - ( 60'd1 << 55 ) : r ;
         r = b [ 50 ] ? r - ( 60'd1 << 54 ) : r ;
         r = b [ 49 ] ? r - ( 60'd1 << 53 ) : r ;
         r = b [ 48 ] ? r - ( 60'd1 << 52 ) : r ;
         r = b [ 47 ] ? r - ( 60'd1 << 51 ) : r ;
         r = b [ 46 ] ? r - ( 60'd1 << 50 ) : r ;
         r = b [ 45 ] ? r - ( 60'd1 << 49 ) : r ;
         r = b [ 44 ] ? r - ( 60'd1 << 48 ) : r ;
         r = b [ 43 ] ? r - ( 60'd1 << 47 ) : r ;
         r = b [ 42 ] ? r - ( 60'd1 << 46 ) : r ;
         r = b [ 41 ] ? r - ( 60'd1 << 45 ) : r ;
         r = b [ 40 ] ? r - ( 60'd1 << 44 ) : r ;
         r = b [ 39 ] ? r - ( 60'd1 << 43 ) : r ;
         r = b [ 38 ] ? r - ( 60'd1 << 42 ) : r ;
         r = b [ 37 ] ? r - ( 60'd1 << 41 ) : r ;
         r = b [ 36 ] ? r - ( 60'd1 << 40 ) : r ;
         r = b [ 35 ] ? r - ( 60'd1 << 39 ) : r ;
         r = b [ 34 ] ? r - ( 60'd1 << 38 ) : r ;
         r = b [ 33 ] ? r - ( 60'd1 << 37 ) : r ;
         r = b [ 32 ] ? r - ( 60'd1 << 36 ) : r ;
         r = b [ 31 ] ? r - ( 60'd1 << 35 ) : r ;
         r = b [ 30 ] ? r - ( 60'd1 << 34 ) : r ;
         r = b [ 29 ] ? r - ( 60'd1 << 33 ) : r ;
         r = b [ 28 ] ? r - ( 60'd1 << 32 ) : r ;
         r = b [ 27 ] ? r - ( 60'd1 << 31 ) : r ;
         r = b [ 26 ] ? r - ( 60'd1 << 30 ) : r ;
         r = b [ 25 ] ? r - ( 60'd1 << 29 ) : r ;
         r = b [ 24 ] ? r - ( 60'd1 << 28 ) : r ;
         r = b [ 23 ] ? r - ( 60'd1 << 27 ) : r ;
         r = b [ 22 ] ? r - ( 60'd1 << 26 ) : r ;
         r = b [ 21 ] ? r - ( 60'd1 << 25 ) : r ;
         r = b [ 20 ] ? r - ( 60'd1 << 24 ) : r ;
         r = b [ 19 ] ? r - ( 60'd1 << 23 ) : r ;
         r = b [ 18 ] ? r - ( 60'd1 << 22 ) : r ;
         r = b [ 17 ] ? r - ( 60'd1 << 21 ) : r ;
         r = b [ 16 ] ? r - ( 60'd1 << 20 ) : r ;
         r = b [ 15 ] ? r - ( 60'd1 << 19 ) : r ;
         r = b [ 14 ] ? r - ( 60'd1 << 18 ) : r ;
         r = b [ 13 ] ? r - ( 60'd1 << 17 ) : r ;
         r = b [ 12 ] ? r - ( 60'd1 << 16 ) : r ;
         r = b [ 11 ] ? r - ( 60'd1 << 15 ) : r ;
         r = b [ 10 ] ? r - ( 60'd1 << 14 ) : r ;
         r = b [ 9 ] ? r - ( 60'd1 << 13 ) : r ;
         r = b [ 8 ] ? r - ( 60'd1 << 12 ) : r ;
         r = b [ 7 ] ? r - ( 60'd1 << 11 ) : r ;
         r = b [ 6 ] ? r - ( 60'd1 << 10 ) : r ;
         r = b [ 5 ] ? r - ( 60'd1 << 9 ) : r ;
         r = b [ 4 ] ? r - ( 60'd1 << 8 ) : r ;
         r = b [ 3 ] ? r - ( 60'd1 << 7 ) : r ;
         r = b [ 2 ] ? r - ( 60'd1 << 6 ) : r ;
         r = b [ 1 ] ? r - ( 60'd1 << 5 ) : r ;
         r = b [ 0 ] ? r - ( 60'd1 << 4 ) : r ;
      end

// Bit by Bit Multiply & Divide + Modulus
// Copyright © 2022 by Gregory Scott Callen
// All Rights Reserved.

      if (( b << 3n ) <= r ) begin
         n = n | 60'd8;
         r = b [ 56 ] ? r - ( 60'd1 << 59 ) : r ;
         r = b [ 55 ] ? r - ( 60'd1 << 58 ) : r ;
         r = b [ 54 ] ? r - ( 60'd1 << 57 ) : r ;
         r = b [ 53 ] ? r - ( 60'd1 << 56 ) : r ;
         r = b [ 52 ] ? r - ( 60'd1 << 55 ) : r ;
         r = b [ 51 ] ? r - ( 60'd1 << 54 ) : r ;
         r = b [ 50 ] ? r - ( 60'd1 << 53 ) : r ;
         r = b [ 49 ] ? r - ( 60'd1 << 52 ) : r ;
         r = b [ 48 ] ? r - ( 60'd1 << 51 ) : r ;
         r = b [ 47 ] ? r - ( 60'd1 << 50 ) : r ;
         r = b [ 46 ] ? r - ( 60'd1 << 49 ) : r ;
         r = b [ 45 ] ? r - ( 60'd1 << 48 ) : r ;
         r = b [ 44 ] ? r - ( 60'd1 << 47 ) : r ;
         r = b [ 43 ] ? r - ( 60'd1 << 46 ) : r ;
         r = b [ 42 ] ? r - ( 60'd1 << 45 ) : r ;
         r = b [ 41 ] ? r - ( 60'd1 << 44 ) : r ;
         r = b [ 40 ] ? r - ( 60'd1 << 43 ) : r ;
         r = b [ 39 ] ? r - ( 60'd1 << 42 ) : r ;
         r = b [ 38 ] ? r - ( 60'd1 << 41 ) : r ;
         r = b [ 37 ] ? r - ( 60'd1 << 40 ) : r ;
         r = b [ 36 ] ? r - ( 60'd1 << 39 ) : r ;
         r = b [ 35 ] ? r - ( 60'd1 << 38 ) : r ;
         r = b [ 34 ] ? r - ( 60'd1 << 37 ) : r ;
         r = b [ 33 ] ? r - ( 60'd1 << 36 ) : r ;
         r = b [ 32 ] ? r - ( 60'd1 << 35 ) : r ;
         r = b [ 31 ] ? r - ( 60'd1 << 34 ) : r ;
         r = b [ 30 ] ? r - ( 60'd1 << 33 ) : r ;
         r = b [ 29 ] ? r - ( 60'd1 << 32 ) : r ;
         r = b [ 28 ] ? r - ( 60'd1 << 31 ) : r ;
         r = b [ 27 ] ? r - ( 60'd1 << 30 ) : r ;
         r = b [ 26 ] ? r - ( 60'd1 << 29 ) : r ;
         r = b [ 25 ] ? r - ( 60'd1 << 28 ) : r ;
         r = b [ 24 ] ? r - ( 60'd1 << 27 ) : r ;
         r = b [ 23 ] ? r - ( 60'd1 << 26 ) : r ;
         r = b [ 22 ] ? r - ( 60'd1 << 25 ) : r ;
         r = b [ 21 ] ? r - ( 60'd1 << 24 ) : r ;
         r = b [ 20 ] ? r - ( 60'd1 << 23 ) : r ;
         r = b [ 19 ] ? r - ( 60'd1 << 22 ) : r ;
         r = b [ 18 ] ? r - ( 60'd1 << 21 ) : r ;
         r = b [ 17 ] ? r - ( 60'd1 << 20 ) : r ;
         r = b [ 16 ] ? r - ( 60'd1 << 19 ) : r ;
         r = b [ 15 ] ? r - ( 60'd1 << 18 ) : r ;
         r = b [ 14 ] ? r - ( 60'd1 << 17 ) : r ;
         r = b [ 13 ] ? r - ( 60'd1 << 16 ) : r ;
         r = b [ 12 ] ? r - ( 60'd1 << 15 ) : r ;
         r = b [ 11 ] ? r - ( 60'd1 << 14 ) : r ;
         r = b [ 10 ] ? r - ( 60'd1 << 13 ) : r ;
         r = b [ 9 ] ? r - ( 60'd1 << 12 ) : r ;
         r = b [ 8 ] ? r - ( 60'd1 << 11 ) : r ;
         r = b [ 7 ] ? r - ( 60'd1 << 10 ) : r ;
         r = b [ 6 ] ? r - ( 60'd1 << 9 ) : r ;
         r = b [ 5 ] ? r - ( 60'd1 << 8 ) : r ;
         r = b [ 4 ] ? r - ( 60'd1 << 7 ) : r ;
         r = b [ 3 ] ? r - ( 60'd1 << 6 ) : r ;
         r = b [ 2 ] ? r - ( 60'd1 << 5 ) : r ;
         r = b [ 1 ] ? r - ( 60'd1 << 4 ) : r ;
         r = b [ 0 ] ? r - ( 60'd1 << 3 ) : r ;
      end

// Bit by Bit Multiply & Divide + Modulus
// Copyright © 2022 by Gregory Scott Callen
// All Rights Reserved.

      if (( b << 2n ) <= r ) begin
         n = n | 60'd4;
         r = b [ 57 ] ? r - ( 60'd1 << 59 ) : r ;
         r = b [ 56 ] ? r - ( 60'd1 << 58 ) : r ;
         r = b [ 55 ] ? r - ( 60'd1 << 57 ) : r ;
         r = b [ 54 ] ? r - ( 60'd1 << 56 ) : r ;
         r = b [ 53 ] ? r - ( 60'd1 << 55 ) : r ;
         r = b [ 52 ] ? r - ( 60'd1 << 54 ) : r ;
         r = b [ 51 ] ? r - ( 60'd1 << 53 ) : r ;
         r = b [ 50 ] ? r - ( 60'd1 << 52 ) : r ;
         r = b [ 49 ] ? r - ( 60'd1 << 51 ) : r ;
         r = b [ 48 ] ? r - ( 60'd1 << 50 ) : r ;
         r = b [ 47 ] ? r - ( 60'd1 << 49 ) : r ;
         r = b [ 46 ] ? r - ( 60'd1 << 48 ) : r ;
         r = b [ 45 ] ? r - ( 60'd1 << 47 ) : r ;
         r = b [ 44 ] ? r - ( 60'd1 << 46 ) : r ;
         r = b [ 43 ] ? r - ( 60'd1 << 45 ) : r ;
         r = b [ 42 ] ? r - ( 60'd1 << 44 ) : r ;
         r = b [ 41 ] ? r - ( 60'd1 << 43 ) : r ;
         r = b [ 40 ] ? r - ( 60'd1 << 42 ) : r ;
         r = b [ 39 ] ? r - ( 60'd1 << 41 ) : r ;
         r = b [ 38 ] ? r - ( 60'd1 << 40 ) : r ;
         r = b [ 37 ] ? r - ( 60'd1 << 39 ) : r ;
         r = b [ 36 ] ? r - ( 60'd1 << 38 ) : r ;
         r = b [ 35 ] ? r - ( 60'd1 << 37 ) : r ;
         r = b [ 34 ] ? r - ( 60'd1 << 36 ) : r ;
         r = b [ 33 ] ? r - ( 60'd1 << 35 ) : r ;
         r = b [ 32 ] ? r - ( 60'd1 << 34 ) : r ;
         r = b [ 31 ] ? r - ( 60'd1 << 33 ) : r ;
         r = b [ 30 ] ? r - ( 60'd1 << 32 ) : r ;
         r = b [ 29 ] ? r - ( 60'd1 << 31 ) : r ;
         r = b [ 28 ] ? r - ( 60'd1 << 30 ) : r ;
         r = b [ 27 ] ? r - ( 60'd1 << 29 ) : r ;
         r = b [ 26 ] ? r - ( 60'd1 << 28 ) : r ;
         r = b [ 25 ] ? r - ( 60'd1 << 27 ) : r ;
         r = b [ 24 ] ? r - ( 60'd1 << 26 ) : r ;
         r = b [ 23 ] ? r - ( 60'd1 << 25 ) : r ;
         r = b [ 22 ] ? r - ( 60'd1 << 24 ) : r ;
         r = b [ 21 ] ? r - ( 60'd1 << 23 ) : r ;
         r = b [ 20 ] ? r - ( 60'd1 << 22 ) : r ;
         r = b [ 19 ] ? r - ( 60'd1 << 21 ) : r ;
         r = b [ 18 ] ? r - ( 60'd1 << 20 ) : r ;
         r = b [ 17 ] ? r - ( 60'd1 << 19 ) : r ;
         r = b [ 16 ] ? r - ( 60'd1 << 18 ) : r ;
         r = b [ 15 ] ? r - ( 60'd1 << 17 ) : r ;
         r = b [ 14 ] ? r - ( 60'd1 << 16 ) : r ;
         r = b [ 13 ] ? r - ( 60'd1 << 15 ) : r ;
         r = b [ 12 ] ? r - ( 60'd1 << 14 ) : r ;
         r = b [ 11 ] ? r - ( 60'd1 << 13 ) : r ;
         r = b [ 10 ] ? r - ( 60'd1 << 12 ) : r ;
         r = b [ 9 ] ? r - ( 60'd1 << 11 ) : r ;
         r = b [ 8 ] ? r - ( 60'd1 << 10 ) : r ;
         r = b [ 7 ] ? r - ( 60'd1 << 9 ) : r ;
         r = b [ 6 ] ? r - ( 60'd1 << 8 ) : r ;
         r = b [ 5 ] ? r - ( 60'd1 << 7 ) : r ;
         r = b [ 4 ] ? r - ( 60'd1 << 6 ) : r ;
         r = b [ 3 ] ? r - ( 60'd1 << 5 ) : r ;
         r = b [ 2 ] ? r - ( 60'd1 << 4 ) : r ;
         r = b [ 1 ] ? r - ( 60'd1 << 3 ) : r ;
         r = b [ 0 ] ? r - ( 60'd1 << 2 ) : r ;
      end

// Bit by Bit Multiply & Divide + Modulus
// Copyright © 2022 by Gregory Scott Callen
// All Rights Reserved.

      if (( b << 1n ) <= r ) begin
         n = n | 60'd2;
         r = b [ 58 ] ? r - ( 60'd1 << 59 ) : r ;
         r = b [ 57 ] ? r - ( 60'd1 << 58 ) : r ;
         r = b [ 56 ] ? r - ( 60'd1 << 57 ) : r ;
         r = b [ 55 ] ? r - ( 60'd1 << 56 ) : r ;
         r = b [ 54 ] ? r - ( 60'd1 << 55 ) : r ;
         r = b [ 53 ] ? r - ( 60'd1 << 54 ) : r ;
         r = b [ 52 ] ? r - ( 60'd1 << 53 ) : r ;
         r = b [ 51 ] ? r - ( 60'd1 << 52 ) : r ;
         r = b [ 50 ] ? r - ( 60'd1 << 51 ) : r ;
         r = b [ 49 ] ? r - ( 60'd1 << 50 ) : r ;
         r = b [ 48 ] ? r - ( 60'd1 << 49 ) : r ;
         r = b [ 47 ] ? r - ( 60'd1 << 48 ) : r ;
         r = b [ 46 ] ? r - ( 60'd1 << 47 ) : r ;
         r = b [ 45 ] ? r - ( 60'd1 << 46 ) : r ;
         r = b [ 44 ] ? r - ( 60'd1 << 45 ) : r ;
         r = b [ 43 ] ? r - ( 60'd1 << 44 ) : r ;
         r = b [ 42 ] ? r - ( 60'd1 << 43 ) : r ;
         r = b [ 41 ] ? r - ( 60'd1 << 42 ) : r ;
         r = b [ 40 ] ? r - ( 60'd1 << 41 ) : r ;
         r = b [ 39 ] ? r - ( 60'd1 << 40 ) : r ;
         r = b [ 38 ] ? r - ( 60'd1 << 39 ) : r ;
         r = b [ 37 ] ? r - ( 60'd1 << 38 ) : r ;
         r = b [ 36 ] ? r - ( 60'd1 << 37 ) : r ;
         r = b [ 35 ] ? r - ( 60'd1 << 36 ) : r ;
         r = b [ 34 ] ? r - ( 60'd1 << 35 ) : r ;
         r = b [ 33 ] ? r - ( 60'd1 << 34 ) : r ;
         r = b [ 32 ] ? r - ( 60'd1 << 33 ) : r ;
         r = b [ 31 ] ? r - ( 60'd1 << 32 ) : r ;
         r = b [ 30 ] ? r - ( 60'd1 << 31 ) : r ;
         r = b [ 29 ] ? r - ( 60'd1 << 30 ) : r ;
         r = b [ 28 ] ? r - ( 60'd1 << 29 ) : r ;
         r = b [ 27 ] ? r - ( 60'd1 << 28 ) : r ;
         r = b [ 26 ] ? r - ( 60'd1 << 27 ) : r ;
         r = b [ 25 ] ? r - ( 60'd1 << 26 ) : r ;
         r = b [ 24 ] ? r - ( 60'd1 << 25 ) : r ;
         r = b [ 23 ] ? r - ( 60'd1 << 24 ) : r ;
         r = b [ 22 ] ? r - ( 60'd1 << 23 ) : r ;
         r = b [ 21 ] ? r - ( 60'd1 << 22 ) : r ;
         r = b [ 20 ] ? r - ( 60'd1 << 21 ) : r ;
         r = b [ 19 ] ? r - ( 60'd1 << 20 ) : r ;
         r = b [ 18 ] ? r - ( 60'd1 << 19 ) : r ;
         r = b [ 17 ] ? r - ( 60'd1 << 18 ) : r ;
         r = b [ 16 ] ? r - ( 60'd1 << 17 ) : r ;
         r = b [ 15 ] ? r - ( 60'd1 << 16 ) : r ;
         r = b [ 14 ] ? r - ( 60'd1 << 15 ) : r ;
         r = b [ 13 ] ? r - ( 60'd1 << 14 ) : r ;
         r = b [ 12 ] ? r - ( 60'd1 << 13 ) : r ;
         r = b [ 11 ] ? r - ( 60'd1 << 12 ) : r ;
         r = b [ 10 ] ? r - ( 60'd1 << 11 ) : r ;
         r = b [ 9 ] ? r - ( 60'd1 << 10 ) : r ;
         r = b [ 8 ] ? r - ( 60'd1 << 9 ) : r ;
         r = b [ 7 ] ? r - ( 60'd1 << 8 ) : r ;
         r = b [ 6 ] ? r - ( 60'd1 << 7 ) : r ;
         r = b [ 5 ] ? r - ( 60'd1 << 6 ) : r ;
         r = b [ 4 ] ? r - ( 60'd1 << 5 ) : r ;
         r = b [ 3 ] ? r - ( 60'd1 << 4 ) : r ;
         r = b [ 2 ] ? r - ( 60'd1 << 3 ) : r ;
         r = b [ 1 ] ? r - ( 60'd1 << 2 ) : r ;
         r = b [ 0 ] ? r - ( 60'd1 << 1 ) : r ;
      end

// Bit by Bit Multiply & Divide + Modulus
// Copyright © 2022 by Gregory Scott Callen
// All Rights Reserved.

      if (( b << 0n ) <= r ) begin
         n = n | 60'd1;
         r = b [ 59 ] ? r - ( 60'd1 << 59 ) : r ;
         r = b [ 58 ] ? r - ( 60'd1 << 58 ) : r ;
         r = b [ 57 ] ? r - ( 60'd1 << 57 ) : r ;
         r = b [ 56 ] ? r - ( 60'd1 << 56 ) : r ;
         r = b [ 55 ] ? r - ( 60'd1 << 55 ) : r ;
         r = b [ 54 ] ? r - ( 60'd1 << 54 ) : r ;
         r = b [ 53 ] ? r - ( 60'd1 << 53 ) : r ;
         r = b [ 52 ] ? r - ( 60'd1 << 52 ) : r ;
         r = b [ 51 ] ? r - ( 60'd1 << 51 ) : r ;
         r = b [ 50 ] ? r - ( 60'd1 << 50 ) : r ;
         r = b [ 49 ] ? r - ( 60'd1 << 49 ) : r ;
         r = b [ 48 ] ? r - ( 60'd1 << 48 ) : r ;
         r = b [ 47 ] ? r - ( 60'd1 << 47 ) : r ;
         r = b [ 46 ] ? r - ( 60'd1 << 46 ) : r ;
         r = b [ 45 ] ? r - ( 60'd1 << 45 ) : r ;
         r = b [ 44 ] ? r - ( 60'd1 << 44 ) : r ;
         r = b [ 43 ] ? r - ( 60'd1 << 43 ) : r ;
         r = b [ 42 ] ? r - ( 60'd1 << 42 ) : r ;
         r = b [ 41 ] ? r - ( 60'd1 << 41 ) : r ;
         r = b [ 40 ] ? r - ( 60'd1 << 40 ) : r ;
         r = b [ 39 ] ? r - ( 60'd1 << 39 ) : r ;
         r = b [ 38 ] ? r - ( 60'd1 << 38 ) : r ;
         r = b [ 37 ] ? r - ( 60'd1 << 37 ) : r ;
         r = b [ 36 ] ? r - ( 60'd1 << 36 ) : r ;
         r = b [ 35 ] ? r - ( 60'd1 << 35 ) : r ;
         r = b [ 34 ] ? r - ( 60'd1 << 34 ) : r ;
         r = b [ 33 ] ? r - ( 60'd1 << 33 ) : r ;
         r = b [ 32 ] ? r - ( 60'd1 << 32 ) : r ;
         r = b [ 31 ] ? r - ( 60'd1 << 31 ) : r ;
         r = b [ 30 ] ? r - ( 60'd1 << 30 ) : r ;
         r = b [ 29 ] ? r - ( 60'd1 << 29 ) : r ;
         r = b [ 28 ] ? r - ( 60'd1 << 28 ) : r ;
         r = b [ 27 ] ? r - ( 60'd1 << 27 ) : r ;
         r = b [ 26 ] ? r - ( 60'd1 << 26 ) : r ;
         r = b [ 25 ] ? r - ( 60'd1 << 25 ) : r ;
         r = b [ 24 ] ? r - ( 60'd1 << 24 ) : r ;
         r = b [ 23 ] ? r - ( 60'd1 << 23 ) : r ;
         r = b [ 22 ] ? r - ( 60'd1 << 22 ) : r ;
         r = b [ 21 ] ? r - ( 60'd1 << 21 ) : r ;
         r = b [ 20 ] ? r - ( 60'd1 << 20 ) : r ;
         r = b [ 19 ] ? r - ( 60'd1 << 19 ) : r ;
         r = b [ 18 ] ? r - ( 60'd1 << 18 ) : r ;
         r = b [ 17 ] ? r - ( 60'd1 << 17 ) : r ;
         r = b [ 16 ] ? r - ( 60'd1 << 16 ) : r ;
         r = b [ 15 ] ? r - ( 60'd1 << 15 ) : r ;
         r = b [ 14 ] ? r - ( 60'd1 << 14 ) : r ;
         r = b [ 13 ] ? r - ( 60'd1 << 13 ) : r ;
         r = b [ 12 ] ? r - ( 60'd1 << 12 ) : r ;
         r = b [ 11 ] ? r - ( 60'd1 << 11 ) : r ;
         r = b [ 10 ] ? r - ( 60'd1 << 10 ) : r ;
         r = b [ 9 ] ? r - ( 60'd1 << 9 ) : r ;
         r = b [ 8 ] ? r - ( 60'd1 << 8 ) : r ;
         r = b [ 7 ] ? r - ( 60'd1 << 7 ) : r ;
         r = b [ 6 ] ? r - ( 60'd1 << 6 ) : r ;
         r = b [ 5 ] ? r - ( 60'd1 << 5 ) : r ;
         r = b [ 4 ] ? r - ( 60'd1 << 4 ) : r ;
         r = b [ 3 ] ? r - ( 60'd1 << 3 ) : r ;
         r = b [ 2 ] ? r - ( 60'd1 << 2 ) : r ;
         r = b [ 1 ] ? r - ( 60'd1 << 1 ) : r ;
         r = b [ 0 ] ? r - ( 60'd1 << 0 ) : r ;
      end

// Bit by Bit Multiply & Divide + Modulus
// Copyright © 2022 by Gregory Scott Callen
// All Rights Reserved.

   end

   // 141041 = 90198117197 / 639514 r 423123

endmodule
